// Benchmark "iscas85-original/c3540" written by ABC on Sat Nov 18 15:15:44 2023

module c3540  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  wire new_n73, new_n74, new_n75, new_n77, new_n78, new_n79, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n104, new_n105,
    new_n106, new_n107, new_n108, new_n109, new_n110, new_n111, new_n112,
    new_n113, new_n115, new_n116, new_n117, new_n118, new_n119, new_n120,
    new_n121, new_n123, new_n124, new_n125, new_n126, new_n127, new_n128,
    new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n277, new_n278,
    new_n279, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n521, new_n522, new_n523, new_n525, new_n526, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535;
  INV_X1    g000(.A(G8), .ZN(new_n73));
  INV_X1    g001(.A(G9), .ZN(new_n74));
  NAND2_X1  g002(.A1(new_n73), .A2(new_n74), .ZN(new_n75));
  NOR3_X1   g003(.A1(G7), .A2(new_n75), .A3(G10), .ZN(G3519));
  INV_X1    g004(.A(G12), .ZN(new_n77));
  INV_X1    g005(.A(G13), .ZN(new_n78));
  NAND2_X1  g006(.A1(new_n77), .A2(new_n78), .ZN(new_n79));
  NAND2_X1  g007(.A1(G11), .A2(new_n79), .ZN(G3520));
  INV_X1    g008(.A(G3), .ZN(new_n81));
  INV_X1    g009(.A(G2), .ZN(new_n82));
  NOR2_X1   g010(.A1(G1), .A2(new_n82), .ZN(new_n83));
  NAND2_X1  g011(.A1(new_n81), .A2(new_n83), .ZN(new_n84));
  INV_X1    g012(.A(G1), .ZN(new_n85));
  NAND2_X1  g013(.A1(new_n85), .A2(new_n82), .ZN(new_n86));
  OR2_X1    g014(.A1(G3), .A2(new_n86), .ZN(new_n87));
  INV_X1    g015(.A(G7), .ZN(new_n88));
  INV_X1    g016(.A(G11), .ZN(new_n89));
  AOI22_X1  g017(.A1(new_n88), .A2(G30), .B1(new_n89), .B2(G34), .ZN(new_n90));
  INV_X1    g018(.A(G36), .ZN(new_n91));
  INV_X1    g019(.A(G32), .ZN(new_n92));
  OAI221_X1 g020(.A(new_n90), .B1(G13), .B2(new_n91), .C1(G9), .C2(new_n92), .ZN(new_n93));
  INV_X1    g021(.A(G10), .ZN(new_n94));
  AOI22_X1  g022(.A1(new_n94), .A2(G33), .B1(new_n73), .B2(G31), .ZN(new_n95));
  INV_X1    g023(.A(G37), .ZN(new_n96));
  INV_X1    g024(.A(G35), .ZN(new_n97));
  OAI221_X1 g025(.A(new_n95), .B1(G14), .B2(new_n96), .C1(G12), .C2(new_n97), .ZN(new_n98));
  OAI211_X1 g026(.A(new_n84), .B(new_n87), .C1(new_n93), .C2(new_n98), .ZN(new_n99));
  NAND2_X1  g027(.A1(new_n88), .A2(new_n75), .ZN(new_n100));
  OAI21_X1  g028(.A(G34), .B1(G35), .B2(G36), .ZN(new_n101));
  OAI221_X1 g029(.A(new_n99), .B1(new_n84), .B2(new_n100), .C1(new_n87), .C2(new_n101), .ZN(new_n102));
  INV_X1    g030(.A(new_n102), .ZN(G3521));
  INV_X1    g031(.A(G34), .ZN(new_n104));
  OAI22_X1  g032(.A1(new_n104), .A2(G35), .B1(G34), .B2(new_n97), .ZN(new_n105));
  OAI22_X1  g033(.A1(G36), .A2(G37), .B1(new_n91), .B2(new_n96), .ZN(new_n106));
  INV_X1    g034(.A(G33), .ZN(new_n107));
  OAI22_X1  g035(.A1(G32), .A2(G33), .B1(new_n92), .B2(new_n107), .ZN(new_n108));
  INV_X1    g036(.A(G30), .ZN(new_n109));
  INV_X1    g037(.A(G31), .ZN(new_n110));
  OAI22_X1  g038(.A1(new_n109), .A2(G31), .B1(G30), .B2(new_n110), .ZN(new_n111));
  XOR2_X1   g039(.A(new_n108), .B(new_n111), .Z(new_n112));
  XNOR2_X1  g040(.A(new_n106), .B(new_n112), .ZN(new_n113));
  XNOR2_X1  g041(.A(new_n105), .B(new_n113), .ZN(G3522));
  OAI22_X1  g042(.A1(new_n89), .A2(G12), .B1(G11), .B2(new_n77), .ZN(new_n115));
  INV_X1    g043(.A(G14), .ZN(new_n116));
  OAI22_X1  g044(.A1(G13), .A2(G14), .B1(new_n78), .B2(new_n116), .ZN(new_n117));
  OAI22_X1  g045(.A1(G9), .A2(new_n94), .B1(new_n74), .B2(G10), .ZN(new_n118));
  OAI22_X1  g046(.A1(new_n88), .A2(G8), .B1(G7), .B2(new_n73), .ZN(new_n119));
  XOR2_X1   g047(.A(new_n118), .B(new_n119), .Z(new_n120));
  XNOR2_X1  g048(.A(new_n117), .B(new_n120), .ZN(new_n121));
  XOR2_X1   g049(.A(new_n115), .B(new_n121), .Z(G3523));
  INV_X1    g050(.A(G4), .ZN(new_n123));
  NOR2_X1   g051(.A1(G1), .A2(new_n123), .ZN(new_n124));
  NOR2_X1   g052(.A1(new_n81), .A2(new_n123), .ZN(new_n125));
  OAI21_X1  g053(.A(G1), .B1(G2), .B2(new_n125), .ZN(new_n126));
  INV_X1    g054(.A(new_n126), .ZN(new_n127));
  INV_X1    g055(.A(new_n83), .ZN(new_n128));
  NOR2_X1   g056(.A1(new_n81), .A2(new_n128), .ZN(new_n129));
  NOR2_X1   g057(.A1(new_n127), .A2(new_n129), .ZN(new_n130));
  INV_X1    g058(.A(new_n130), .ZN(new_n131));
  NOR3_X1   g059(.A1(new_n78), .A2(new_n124), .A3(new_n131), .ZN(new_n132));
  NAND2_X1  g060(.A1(G3), .A2(new_n78), .ZN(new_n133));
  NAND2_X1  g061(.A1(new_n81), .A2(G4), .ZN(new_n134));
  NAND2_X1  g062(.A1(new_n81), .A2(new_n123), .ZN(new_n135));
  OAI221_X1 g063(.A(new_n133), .B1(new_n116), .B2(new_n134), .C1(G11), .C2(new_n135), .ZN(new_n136));
  AOI221_X1 g064(.A(new_n132), .B1(new_n78), .B2(new_n129), .C1(new_n127), .C2(new_n136), .ZN(new_n137));
  NOR2_X1   g065(.A1(G25), .A2(G26), .ZN(new_n138));
  INV_X1    g066(.A(G6), .ZN(new_n139));
  NAND2_X1  g067(.A1(new_n85), .A2(new_n139), .ZN(new_n140));
  INV_X1    g068(.A(G38), .ZN(new_n141));
  INV_X1    g069(.A(G5), .ZN(new_n142));
  NOR2_X1   g070(.A1(new_n123), .A2(new_n142), .ZN(new_n143));
  NOR3_X1   g071(.A1(new_n85), .A2(new_n82), .A3(new_n143), .ZN(new_n144));
  NOR4_X1   g072(.A1(G5), .A2(new_n140), .A3(new_n141), .A4(new_n144), .ZN(new_n145));
  INV_X1    g073(.A(new_n145), .ZN(new_n146));
  NOR2_X1   g074(.A1(G5), .A2(new_n140), .ZN(new_n147));
  NOR2_X1   g075(.A1(new_n91), .A2(new_n147), .ZN(new_n148));
  INV_X1    g076(.A(G40), .ZN(new_n149));
  OAI21_X1  g077(.A(new_n149), .B1(new_n104), .B2(G49), .ZN(new_n150));
  AOI221_X1 g078(.A(new_n148), .B1(G4), .B2(G35), .C1(new_n123), .C2(new_n150), .ZN(new_n151));
  OAI21_X1  g079(.A(new_n146), .B1(new_n144), .B2(new_n151), .ZN(new_n152));
  OAI21_X1  g080(.A(new_n137), .B1(new_n138), .B2(new_n152), .ZN(new_n153));
  NOR2_X1   g081(.A1(G23), .A2(G24), .ZN(new_n154));
  OR2_X1    g082(.A1(new_n152), .A2(new_n154), .ZN(new_n155));
  NOR2_X1   g083(.A1(new_n137), .A2(new_n155), .ZN(new_n156));
  INV_X1    g084(.A(new_n156), .ZN(new_n157));
  NAND2_X1  g085(.A1(new_n153), .A2(new_n157), .ZN(new_n158));
  NOR2_X1   g086(.A1(G11), .A2(new_n79), .ZN(new_n159));
  OAI222_X1 g087(.A1(G12), .A2(new_n134), .B1(G9), .B2(new_n135), .C1(new_n81), .C2(new_n159), .ZN(new_n160));
  NOR2_X1   g088(.A1(new_n89), .A2(new_n124), .ZN(new_n161));
  AOI222_X1 g089(.A1(new_n127), .A2(new_n160), .B1(new_n89), .B2(new_n129), .C1(new_n130), .C2(new_n161), .ZN(new_n162));
  OAI22_X1  g090(.A1(new_n141), .A2(new_n140), .B1(new_n123), .B2(new_n107), .ZN(new_n163));
  OAI21_X1  g091(.A(new_n116), .B1(new_n92), .B2(G49), .ZN(new_n164));
  AOI221_X1 g092(.A(new_n163), .B1(G34), .B2(new_n140), .C1(new_n123), .C2(new_n164), .ZN(new_n165));
  NOR2_X1   g093(.A1(new_n144), .A2(new_n165), .ZN(new_n166));
  OAI21_X1  g094(.A(new_n162), .B1(new_n138), .B2(new_n166), .ZN(new_n167));
  OR2_X1    g095(.A1(new_n154), .A2(new_n166), .ZN(new_n168));
  OAI21_X1  g096(.A(new_n167), .B1(new_n162), .B2(new_n168), .ZN(new_n169));
  AOI221_X1 g097(.A(G3), .B1(new_n123), .B2(new_n77), .C1(G4), .C2(G39), .ZN(new_n170));
  AOI211_X1 g098(.A(new_n126), .B(new_n170), .C1(G3), .C2(new_n116), .ZN(new_n171));
  OAI33_X1  g099(.A1(new_n81), .A2(G14), .A3(new_n128), .B1(new_n116), .B2(new_n124), .B3(new_n131), .ZN(new_n172));
  INV_X1    g100(.A(new_n138), .ZN(new_n173));
  NOR2_X1   g101(.A1(new_n96), .A2(new_n147), .ZN(new_n174));
  INV_X1    g102(.A(G41), .ZN(new_n175));
  OAI21_X1  g103(.A(new_n175), .B1(new_n97), .B2(G49), .ZN(new_n176));
  AOI221_X1 g104(.A(new_n174), .B1(G4), .B2(G36), .C1(new_n123), .C2(new_n176), .ZN(new_n177));
  NOR2_X1   g105(.A1(new_n144), .A2(new_n177), .ZN(new_n178));
  NOR2_X1   g106(.A1(new_n145), .A2(new_n178), .ZN(new_n179));
  AOI211_X1 g107(.A(new_n171), .B(new_n172), .C1(new_n173), .C2(new_n179), .ZN(new_n180));
  NOR2_X1   g108(.A1(new_n171), .A2(new_n172), .ZN(new_n181));
  OAI21_X1  g109(.A(new_n179), .B1(G23), .B2(G24), .ZN(new_n182));
  NOR2_X1   g110(.A1(new_n181), .A2(new_n182), .ZN(new_n183));
  OR2_X1    g111(.A1(new_n180), .A2(new_n183), .ZN(new_n184));
  OAI21_X1  g112(.A(new_n79), .B1(new_n77), .B2(new_n78), .ZN(new_n185));
  OAI222_X1 g113(.A1(new_n94), .A2(new_n135), .B1(new_n78), .B2(new_n134), .C1(new_n81), .C2(new_n185), .ZN(new_n186));
  NOR2_X1   g114(.A1(new_n77), .A2(new_n124), .ZN(new_n187));
  AOI222_X1 g115(.A1(new_n127), .A2(new_n186), .B1(new_n77), .B2(new_n129), .C1(new_n130), .C2(new_n187), .ZN(new_n188));
  NOR2_X1   g116(.A1(new_n97), .A2(new_n147), .ZN(new_n189));
  INV_X1    g117(.A(G39), .ZN(new_n190));
  OAI21_X1  g118(.A(new_n190), .B1(new_n107), .B2(G49), .ZN(new_n191));
  AOI221_X1 g119(.A(new_n189), .B1(G4), .B2(G34), .C1(new_n123), .C2(new_n191), .ZN(new_n192));
  OAI21_X1  g120(.A(new_n146), .B1(new_n144), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g121(.A(new_n188), .B1(new_n138), .B2(new_n193), .ZN(new_n194));
  INV_X1    g122(.A(new_n193), .ZN(new_n195));
  OAI21_X1  g123(.A(new_n195), .B1(G23), .B2(G24), .ZN(new_n196));
  OAI21_X1  g124(.A(new_n194), .B1(new_n188), .B2(new_n196), .ZN(new_n197));
  OR4_X1    g125(.A1(new_n158), .A2(new_n169), .A3(new_n184), .A4(new_n197), .ZN(new_n198));
  INV_X1    g126(.A(G21), .ZN(new_n199));
  NOR2_X1   g127(.A1(G7), .A2(new_n75), .ZN(new_n200));
  OAI222_X1 g128(.A1(new_n199), .A2(new_n135), .B1(G8), .B2(new_n134), .C1(new_n81), .C2(new_n200), .ZN(new_n201));
  NOR2_X1   g129(.A1(G1), .A2(new_n81), .ZN(new_n202));
  NOR2_X1   g130(.A1(new_n88), .A2(new_n202), .ZN(new_n203));
  AOI222_X1 g131(.A1(new_n127), .A2(new_n201), .B1(new_n88), .B2(new_n129), .C1(new_n130), .C2(new_n203), .ZN(new_n204));
  OAI21_X1  g132(.A(new_n85), .B1(G5), .B2(G6), .ZN(new_n205));
  OR3_X1    g133(.A1(new_n141), .A2(new_n144), .A3(new_n205), .ZN(new_n206));
  INV_X1    g134(.A(G29), .ZN(new_n207));
  INV_X1    g135(.A(G49), .ZN(new_n208));
  AOI21_X1  g136(.A(G10), .B1(G28), .B2(new_n208), .ZN(new_n209));
  OAI22_X1  g137(.A1(new_n123), .A2(new_n207), .B1(G4), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g138(.A(new_n210), .B1(G30), .B2(new_n205), .ZN(new_n211));
  OAI21_X1  g139(.A(new_n206), .B1(new_n144), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g140(.A(new_n204), .B1(new_n138), .B2(new_n212), .ZN(new_n213));
  INV_X1    g141(.A(new_n213), .ZN(new_n214));
  NOR3_X1   g142(.A1(new_n154), .A2(new_n212), .A3(new_n204), .ZN(new_n215));
  NOR2_X1   g143(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI222_X1 g144(.A1(G8), .A2(new_n135), .B1(new_n81), .B2(new_n94), .C1(G11), .C2(new_n134), .ZN(new_n217));
  NOR2_X1   g145(.A1(new_n94), .A2(new_n202), .ZN(new_n218));
  AOI222_X1 g146(.A1(new_n127), .A2(new_n217), .B1(new_n94), .B2(new_n129), .C1(new_n130), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g147(.A(new_n78), .B1(new_n110), .B2(G49), .ZN(new_n220));
  AOI222_X1 g148(.A1(G4), .A2(G32), .B1(new_n123), .B2(new_n220), .C1(G33), .C2(new_n205), .ZN(new_n221));
  OAI21_X1  g149(.A(new_n206), .B1(new_n144), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g150(.A(new_n219), .B1(new_n138), .B2(new_n222), .ZN(new_n223));
  INV_X1    g151(.A(G22), .ZN(new_n224));
  OAI21_X1  g152(.A(new_n75), .B1(new_n73), .B2(new_n74), .ZN(new_n225));
  OAI222_X1 g153(.A1(new_n224), .A2(new_n135), .B1(G9), .B2(new_n134), .C1(new_n81), .C2(new_n225), .ZN(new_n226));
  NOR2_X1   g154(.A1(new_n73), .A2(new_n202), .ZN(new_n227));
  AOI222_X1 g155(.A1(new_n127), .A2(new_n226), .B1(new_n73), .B2(new_n129), .C1(new_n130), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g156(.A(new_n89), .B1(new_n207), .B2(G49), .ZN(new_n229));
  AOI222_X1 g157(.A1(G4), .A2(G30), .B1(new_n123), .B2(new_n229), .C1(G31), .C2(new_n205), .ZN(new_n230));
  OAI21_X1  g158(.A(new_n206), .B1(new_n144), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g159(.A(new_n228), .B1(new_n138), .B2(new_n231), .ZN(new_n232));
  INV_X1    g160(.A(new_n232), .ZN(new_n233));
  NOR3_X1   g161(.A1(new_n154), .A2(new_n231), .A3(new_n228), .ZN(new_n234));
  NOR2_X1   g162(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR3_X1   g163(.A1(new_n74), .A2(new_n202), .A3(new_n131), .ZN(new_n236));
  OAI222_X1 g164(.A1(new_n94), .A2(new_n134), .B1(new_n81), .B2(G9), .C1(new_n88), .C2(new_n135), .ZN(new_n237));
  AOI221_X1 g165(.A(new_n236), .B1(new_n74), .B2(new_n129), .C1(new_n127), .C2(new_n237), .ZN(new_n238));
  OAI21_X1  g166(.A(new_n77), .B1(new_n109), .B2(G49), .ZN(new_n239));
  AOI222_X1 g167(.A1(G32), .A2(new_n205), .B1(G4), .B2(G31), .C1(new_n123), .C2(new_n239), .ZN(new_n240));
  OAI21_X1  g168(.A(new_n206), .B1(new_n144), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g169(.A(new_n238), .B1(new_n138), .B2(new_n241), .ZN(new_n242));
  OR3_X1    g170(.A1(new_n154), .A2(new_n241), .A3(new_n238), .ZN(new_n243));
  AND2_X1   g171(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OR3_X1    g172(.A1(new_n154), .A2(new_n222), .A3(new_n219), .ZN(new_n245));
  NAND2_X1  g173(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g174(.A(new_n246), .ZN(new_n247));
  NAND4_X1  g175(.A1(new_n216), .A2(new_n223), .A3(new_n235), .A4(new_n247), .ZN(new_n248));
  NOR2_X1   g176(.A1(new_n198), .A2(new_n248), .ZN(G3524));
  AOI21_X1  g177(.A(new_n234), .B1(new_n242), .B2(new_n246), .ZN(new_n250));
  NOR2_X1   g178(.A1(new_n233), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g179(.A(new_n213), .B1(new_n215), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g180(.A1(new_n162), .A2(new_n168), .ZN(new_n253));
  INV_X1    g181(.A(new_n167), .ZN(new_n254));
  INV_X1    g182(.A(new_n194), .ZN(new_n255));
  NOR2_X1   g183(.A1(new_n188), .A2(new_n196), .ZN(new_n256));
  AOI211_X1 g184(.A(new_n156), .B(new_n256), .C1(new_n153), .C2(new_n183), .ZN(new_n257));
  NOR3_X1   g185(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g186(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g187(.A(new_n252), .B1(new_n248), .B2(new_n259), .ZN(G3525));
  INV_X1    g188(.A(G47), .ZN(new_n261));
  INV_X1    g189(.A(G48), .ZN(new_n262));
  INV_X1    g190(.A(G27), .ZN(new_n263));
  NOR2_X1   g191(.A1(new_n263), .A2(new_n87), .ZN(new_n264));
  INV_X1    g192(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g193(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g194(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g195(.A1(new_n181), .A2(new_n267), .ZN(new_n268));
  OAI33_X1  g196(.A1(new_n180), .A2(new_n183), .A3(new_n268), .B1(new_n181), .B2(new_n267), .B3(new_n182), .ZN(new_n269));
  NOR2_X1   g197(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g198(.A1(new_n183), .A2(new_n267), .ZN(new_n271));
  NOR2_X1   g199(.A1(new_n137), .A2(new_n267), .ZN(new_n272));
  INV_X1    g200(.A(new_n272), .ZN(new_n273));
  OAI22_X1  g201(.A1(new_n158), .A2(new_n272), .B1(new_n155), .B2(new_n273), .ZN(new_n274));
  XOR2_X1   g202(.A(new_n271), .B(new_n274), .Z(new_n275));
  NOR3_X1   g203(.A1(new_n270), .A2(new_n275), .A3(new_n261), .ZN(G3526));
  NOR2_X1   g204(.A1(new_n142), .A2(new_n87), .ZN(new_n277));
  NOR2_X1   g205(.A1(new_n259), .A2(new_n266), .ZN(new_n278));
  INV_X1    g206(.A(new_n278), .ZN(new_n279));
  OAI22_X1  g207(.A1(new_n100), .A2(new_n277), .B1(G1), .B2(new_n279), .ZN(G3527));
  INV_X1    g208(.A(new_n277), .ZN(new_n281));
  NAND2_X1  g209(.A1(new_n82), .A2(new_n81), .ZN(new_n282));
  OAI21_X1  g210(.A(new_n85), .B1(new_n139), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g211(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AOI211_X1 g212(.A(new_n270), .B(new_n284), .C1(new_n261), .C2(new_n269), .ZN(new_n285));
  OAI21_X1  g213(.A(new_n83), .B1(new_n81), .B2(G23), .ZN(new_n286));
  INV_X1    g214(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g215(.A1(new_n86), .A2(new_n135), .ZN(new_n288));
  NAND3_X1  g216(.A1(new_n88), .A2(new_n75), .A3(G6), .ZN(new_n289));
  OAI21_X1  g217(.A(new_n289), .B1(G6), .B2(new_n120), .ZN(new_n290));
  NAND4_X1  g218(.A1(G11), .A2(new_n79), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  OAI211_X1 g219(.A(new_n287), .B(new_n291), .C1(new_n116), .C2(new_n288), .ZN(new_n292));
  NAND2_X1  g220(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  INV_X1    g221(.A(G25), .ZN(new_n294));
  NOR4_X1   g222(.A1(new_n81), .A2(new_n294), .A3(G24), .A4(G26), .ZN(new_n295));
  INV_X1    g223(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g224(.A(new_n296), .B1(G42), .B2(G46), .ZN(new_n297));
  INV_X1    g225(.A(G24), .ZN(new_n298));
  OAI21_X1  g226(.A(G26), .B1(new_n81), .B2(new_n298), .ZN(new_n299));
  NOR3_X1   g227(.A1(new_n81), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  INV_X1    g228(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g229(.A(new_n299), .B1(G3), .B2(G25), .ZN(new_n302));
  INV_X1    g230(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g231(.A1(G43), .A2(new_n301), .B1(G45), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g232(.A(G3), .B1(G24), .B2(new_n173), .ZN(new_n305));
  OAI211_X1 g233(.A(new_n297), .B(new_n304), .C1(new_n149), .C2(new_n305), .ZN(new_n306));
  AOI21_X1  g234(.A(new_n123), .B1(G39), .B2(new_n301), .ZN(new_n307));
  NOR2_X1   g235(.A1(new_n81), .A2(new_n303), .ZN(new_n308));
  INV_X1    g236(.A(G44), .ZN(new_n309));
  INV_X1    g237(.A(new_n305), .ZN(new_n310));
  NOR2_X1   g238(.A1(G26), .A2(new_n310), .ZN(new_n311));
  OAI221_X1 g239(.A(new_n307), .B1(new_n175), .B2(new_n308), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  OAI22_X1  g240(.A1(G9), .A2(new_n300), .B1(G11), .B2(new_n308), .ZN(new_n313));
  NOR2_X1   g241(.A1(new_n94), .A2(G22), .ZN(new_n314));
  OAI21_X1  g242(.A(new_n123), .B1(new_n295), .B2(new_n314), .ZN(new_n315));
  OAI22_X1  g243(.A1(G13), .A2(new_n300), .B1(G7), .B2(new_n302), .ZN(new_n316));
  AOI211_X1 g244(.A(new_n315), .B(new_n316), .C1(new_n77), .C2(new_n310), .ZN(new_n317));
  OAI21_X1  g245(.A(new_n317), .B1(G8), .B2(new_n311), .ZN(new_n318));
  OAI22_X1  g246(.A1(new_n306), .A2(new_n312), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g247(.A1(new_n123), .A2(new_n282), .ZN(new_n320));
  AOI221_X1 g248(.A(new_n293), .B1(new_n286), .B2(new_n319), .C1(new_n269), .C2(new_n320), .ZN(new_n321));
  OR2_X1    g249(.A1(new_n285), .A2(new_n321), .ZN(G3528));
  OAI21_X1  g250(.A(new_n298), .B1(new_n144), .B2(new_n151), .ZN(new_n323));
  OR2_X1    g251(.A1(new_n166), .A2(new_n178), .ZN(new_n324));
  NAND3_X1  g252(.A1(G24), .A2(new_n166), .A3(new_n152), .ZN(new_n325));
  OAI33_X1  g253(.A1(new_n323), .A2(new_n324), .A3(new_n193), .B1(new_n179), .B2(new_n195), .B3(new_n325), .ZN(new_n326));
  INV_X1    g254(.A(new_n326), .ZN(new_n327));
  OAI22_X1  g255(.A1(new_n266), .A2(new_n327), .B1(new_n198), .B2(new_n267), .ZN(new_n328));
  NAND2_X1  g256(.A1(G47), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g257(.A1(new_n245), .A2(new_n266), .ZN(new_n330));
  OAI21_X1  g258(.A(new_n223), .B1(new_n219), .B2(new_n267), .ZN(new_n331));
  AOI21_X1  g259(.A(new_n330), .B1(new_n245), .B2(new_n331), .ZN(new_n332));
  INV_X1    g260(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g261(.A1(new_n278), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g262(.A(new_n334), .B1(new_n278), .B2(new_n333), .ZN(new_n335));
  AOI21_X1  g263(.A(new_n284), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g264(.A(new_n336), .B1(new_n329), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g265(.A1(new_n116), .A2(G42), .ZN(new_n338));
  OAI22_X1  g266(.A1(G12), .A2(new_n305), .B1(new_n295), .B2(new_n338), .ZN(new_n339));
  OAI22_X1  g267(.A1(G11), .A2(new_n300), .B1(new_n175), .B2(new_n302), .ZN(new_n340));
  OAI221_X1 g268(.A(new_n307), .B1(G13), .B2(new_n308), .C1(new_n149), .C2(new_n311), .ZN(new_n341));
  NOR2_X1   g269(.A1(G18), .A2(G22), .ZN(new_n342));
  OAI221_X1 g270(.A(new_n123), .B1(new_n295), .B2(new_n342), .C1(G8), .C2(new_n305), .ZN(new_n343));
  NOR2_X1   g271(.A1(new_n74), .A2(G21), .ZN(new_n344));
  INV_X1    g272(.A(G19), .ZN(new_n345));
  OAI22_X1  g273(.A1(new_n300), .A2(new_n344), .B1(new_n345), .B2(new_n302), .ZN(new_n346));
  INV_X1    g274(.A(G20), .ZN(new_n347));
  OAI22_X1  g275(.A1(new_n347), .A2(new_n311), .B1(G7), .B2(new_n308), .ZN(new_n348));
  OAI33_X1  g276(.A1(new_n339), .A2(new_n340), .A3(new_n341), .B1(new_n343), .B2(new_n346), .B3(new_n348), .ZN(new_n349));
  INV_X1    g277(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g278(.A1(new_n82), .A2(G4), .ZN(new_n351));
  OAI221_X1 g279(.A(new_n284), .B1(new_n287), .B2(new_n350), .C1(new_n333), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g280(.A1(new_n337), .A2(new_n352), .ZN(G3529));
  NAND4_X1  g281(.A1(new_n81), .A2(new_n116), .A3(new_n83), .A4(new_n185), .ZN(new_n354));
  NAND2_X1  g282(.A1(new_n84), .A2(new_n86), .ZN(new_n355));
  OR2_X1    g283(.A1(new_n261), .A2(new_n328), .ZN(new_n356));
  OAI21_X1  g284(.A(new_n244), .B1(new_n238), .B2(new_n267), .ZN(new_n357));
  OAI21_X1  g285(.A(new_n357), .B1(new_n243), .B2(new_n267), .ZN(new_n358));
  OAI21_X1  g286(.A(new_n235), .B1(new_n228), .B2(new_n265), .ZN(new_n359));
  INV_X1    g287(.A(new_n359), .ZN(new_n360));
  OAI22_X1  g288(.A1(new_n234), .A2(new_n360), .B1(new_n264), .B2(new_n360), .ZN(new_n361));
  INV_X1    g289(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g290(.A1(new_n332), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g291(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g292(.A(new_n248), .ZN(new_n365));
  OR2_X1    g293(.A1(new_n365), .A2(new_n328), .ZN(new_n366));
  NOR2_X1   g294(.A1(new_n261), .A2(new_n366), .ZN(new_n367));
  OAI22_X1  g295(.A1(new_n364), .A2(new_n367), .B1(new_n363), .B2(new_n366), .ZN(new_n368));
  INV_X1    g296(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g297(.A(new_n252), .B1(new_n365), .B2(new_n278), .ZN(new_n370));
  NOR2_X1   g298(.A1(new_n264), .A2(new_n360), .ZN(new_n371));
  OAI21_X1  g299(.A(new_n243), .B1(new_n330), .B2(new_n357), .ZN(new_n372));
  OAI22_X1  g300(.A1(new_n234), .A2(new_n360), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g301(.A(new_n370), .B(new_n373), .ZN(new_n374));
  AOI21_X1  g302(.A(new_n355), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g303(.A(new_n375), .B1(new_n369), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g304(.A1(G7), .A2(G10), .ZN(new_n377));
  AOI22_X1  g305(.A1(G7), .A2(new_n74), .B1(new_n225), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g306(.A(new_n354), .B(new_n376), .C1(new_n86), .C2(new_n378), .ZN(G3530));
  INV_X1    g307(.A(new_n284), .ZN(new_n380));
  AOI211_X1 g308(.A(new_n81), .B(G9), .C1(new_n298), .C2(new_n138), .ZN(new_n381));
  NOR2_X1   g309(.A1(new_n88), .A2(G19), .ZN(new_n382));
  OAI21_X1  g310(.A(new_n123), .B1(new_n295), .B2(new_n382), .ZN(new_n383));
  OAI22_X1  g311(.A1(new_n300), .A2(new_n314), .B1(new_n347), .B2(new_n302), .ZN(new_n384));
  NOR3_X1   g312(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI221_X1 g313(.A(new_n385), .B1(G8), .B2(new_n308), .C1(new_n199), .C2(new_n311), .ZN(new_n386));
  AOI21_X1  g314(.A(new_n311), .B1(new_n175), .B2(new_n133), .ZN(new_n387));
  OAI21_X1  g315(.A(new_n296), .B1(G39), .B2(G43), .ZN(new_n388));
  OAI211_X1 g316(.A(G4), .B(new_n388), .C1(G3), .C2(G14), .ZN(new_n389));
  INV_X1    g317(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g318(.A1(new_n77), .A2(G40), .ZN(new_n391));
  OAI221_X1 g319(.A(new_n390), .B1(new_n302), .B2(new_n338), .C1(new_n300), .C2(new_n391), .ZN(new_n392));
  OAI21_X1  g320(.A(new_n386), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g321(.A1(new_n162), .A2(new_n267), .ZN(new_n394));
  OAI33_X1  g322(.A1(new_n254), .A2(new_n253), .A3(new_n394), .B1(new_n162), .B2(new_n267), .B3(new_n168), .ZN(new_n395));
  AOI221_X1 g323(.A(new_n380), .B1(new_n286), .B2(new_n393), .C1(new_n320), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g324(.A1(new_n188), .A2(new_n267), .ZN(new_n397));
  OAI33_X1  g325(.A1(new_n255), .A2(new_n256), .A3(new_n397), .B1(new_n188), .B2(new_n267), .B3(new_n196), .ZN(new_n398));
  INV_X1    g326(.A(new_n398), .ZN(new_n399));
  INV_X1    g327(.A(G3526), .ZN(new_n400));
  OAI22_X1  g328(.A1(new_n271), .A2(new_n274), .B1(new_n157), .B2(new_n266), .ZN(new_n401));
  OAI211_X1 g329(.A(new_n399), .B(new_n400), .C1(new_n256), .C2(new_n401), .ZN(new_n402));
  NOR2_X1   g330(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  INV_X1    g331(.A(new_n283), .ZN(new_n404));
  XOR2_X1   g332(.A(new_n270), .B(new_n275), .Z(new_n405));
  AOI21_X1  g333(.A(new_n277), .B1(new_n278), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g334(.A1(new_n400), .A2(new_n401), .ZN(new_n407));
  XOR2_X1   g335(.A(new_n407), .B(new_n399), .Z(new_n408));
  INV_X1    g336(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g337(.A(new_n406), .B1(new_n279), .B2(new_n409), .ZN(new_n410));
  AOI221_X1 g338(.A(new_n403), .B1(new_n395), .B2(new_n402), .C1(new_n404), .C2(new_n410), .ZN(new_n411));
  OR2_X1    g339(.A1(new_n396), .A2(new_n411), .ZN(G3531));
  INV_X1    g340(.A(new_n112), .ZN(new_n413));
  AOI22_X1  g341(.A1(new_n74), .A2(G10), .B1(G8), .B2(G9), .ZN(new_n414));
  OAI22_X1  g342(.A1(G6), .A2(new_n413), .B1(new_n289), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g343(.A1(new_n116), .A2(new_n159), .A3(new_n288), .A4(new_n415), .ZN(new_n416));
  OAI211_X1 g344(.A(new_n287), .B(new_n416), .C1(new_n78), .C2(new_n288), .ZN(new_n417));
  NAND2_X1  g345(.A1(new_n284), .A2(new_n417), .ZN(new_n418));
  OAI221_X1 g346(.A(G4), .B1(G14), .B2(new_n300), .C1(new_n190), .C2(new_n311), .ZN(new_n419));
  OAI21_X1  g347(.A(new_n419), .B1(new_n116), .B2(new_n134), .ZN(new_n420));
  INV_X1    g348(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g349(.A(new_n296), .B1(G41), .B2(G45), .ZN(new_n422));
  OAI21_X1  g350(.A(new_n422), .B1(new_n309), .B2(new_n302), .ZN(new_n423));
  AOI21_X1  g351(.A(new_n423), .B1(G42), .B2(new_n301), .ZN(new_n424));
  INV_X1    g352(.A(G43), .ZN(new_n425));
  OAI221_X1 g353(.A(new_n424), .B1(new_n425), .B2(new_n311), .C1(new_n149), .C2(new_n308), .ZN(new_n426));
  OAI221_X1 g354(.A(new_n123), .B1(G12), .B2(new_n300), .C1(G10), .C2(new_n308), .ZN(new_n427));
  NOR2_X1   g355(.A1(G8), .A2(new_n300), .ZN(new_n428));
  INV_X1    g356(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g357(.A(new_n429), .B1(new_n295), .B2(new_n344), .ZN(new_n430));
  AOI221_X1 g358(.A(new_n430), .B1(G22), .B2(new_n303), .C1(new_n89), .C2(new_n310), .ZN(new_n431));
  OAI21_X1  g359(.A(new_n431), .B1(G7), .B2(new_n311), .ZN(new_n432));
  OAI22_X1  g360(.A1(new_n421), .A2(new_n426), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  AOI221_X1 g361(.A(new_n418), .B1(new_n286), .B2(new_n433), .C1(new_n274), .C2(new_n320), .ZN(new_n434));
  INV_X1    g362(.A(new_n434), .ZN(new_n435));
  INV_X1    g363(.A(new_n406), .ZN(new_n436));
  NOR2_X1   g364(.A1(new_n278), .A2(new_n405), .ZN(new_n437));
  OAI221_X1 g365(.A(new_n435), .B1(new_n404), .B2(new_n405), .C1(new_n436), .C2(new_n437), .ZN(G3532));
  OAI21_X1  g366(.A(new_n296), .B1(G40), .B2(G44), .ZN(new_n439));
  OAI21_X1  g367(.A(new_n439), .B1(G14), .B2(new_n305), .ZN(new_n440));
  OAI22_X1  g368(.A1(new_n425), .A2(new_n302), .B1(new_n175), .B2(new_n300), .ZN(new_n441));
  AOI21_X1  g369(.A(new_n123), .B1(new_n78), .B2(new_n301), .ZN(new_n442));
  INV_X1    g370(.A(G42), .ZN(new_n443));
  OAI221_X1 g371(.A(new_n442), .B1(new_n190), .B2(new_n308), .C1(new_n443), .C2(new_n311), .ZN(new_n444));
  AOI21_X1  g372(.A(G4), .B1(G20), .B2(new_n296), .ZN(new_n445));
  OAI21_X1  g373(.A(new_n445), .B1(new_n199), .B2(new_n302), .ZN(new_n446));
  NAND2_X1  g374(.A1(new_n94), .A2(new_n310), .ZN(new_n447));
  OAI21_X1  g375(.A(new_n447), .B1(G7), .B2(new_n300), .ZN(new_n448));
  AOI22_X1  g376(.A1(new_n89), .A2(new_n301), .B1(new_n73), .B2(new_n296), .ZN(new_n449));
  OAI221_X1 g377(.A(new_n449), .B1(G9), .B2(new_n308), .C1(new_n224), .C2(new_n311), .ZN(new_n450));
  OAI33_X1  g378(.A1(new_n440), .A2(new_n441), .A3(new_n444), .B1(new_n446), .B2(new_n448), .B3(new_n450), .ZN(new_n451));
  AOI221_X1 g379(.A(new_n380), .B1(new_n286), .B2(new_n451), .C1(new_n320), .C2(new_n398), .ZN(new_n452));
  INV_X1    g380(.A(new_n452), .ZN(new_n453));
  INV_X1    g381(.A(new_n437), .ZN(new_n454));
  OAI221_X1 g382(.A(new_n281), .B1(new_n409), .B2(new_n454), .C1(new_n408), .C2(new_n437), .ZN(new_n455));
  OAI211_X1 g383(.A(new_n453), .B(new_n455), .C1(new_n404), .C2(new_n408), .ZN(G3533));
  INV_X1    g384(.A(G16), .ZN(new_n457));
  INV_X1    g385(.A(G18), .ZN(new_n458));
  OAI221_X1 g386(.A(new_n445), .B1(new_n457), .B2(new_n295), .C1(new_n458), .C2(new_n311), .ZN(new_n459));
  INV_X1    g387(.A(new_n459), .ZN(new_n460));
  OAI22_X1  g388(.A1(new_n300), .A2(new_n382), .B1(new_n224), .B2(new_n305), .ZN(new_n461));
  AOI21_X1  g389(.A(new_n461), .B1(G17), .B2(new_n303), .ZN(new_n462));
  OAI211_X1 g390(.A(new_n460), .B(new_n462), .C1(new_n199), .C2(new_n308), .ZN(new_n463));
  OAI21_X1  g391(.A(new_n447), .B1(new_n295), .B2(new_n391), .ZN(new_n464));
  AOI21_X1  g392(.A(new_n464), .B1(G39), .B2(new_n303), .ZN(new_n465));
  OAI211_X1 g393(.A(new_n442), .B(new_n465), .C1(G14), .C2(new_n311), .ZN(new_n466));
  OAI21_X1  g394(.A(new_n463), .B1(new_n313), .B2(new_n466), .ZN(new_n467));
  INV_X1    g395(.A(new_n467), .ZN(new_n468));
  OAI221_X1 g396(.A(new_n284), .B1(new_n287), .B2(new_n468), .C1(new_n351), .C2(new_n361), .ZN(new_n469));
  INV_X1    g397(.A(new_n358), .ZN(new_n470));
  OR2_X1    g398(.A1(new_n333), .A2(new_n356), .ZN(new_n471));
  OAI21_X1  g399(.A(new_n372), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XOR2_X1   g400(.A(new_n362), .B(new_n472), .Z(new_n473));
  NAND2_X1  g401(.A1(new_n367), .A2(new_n370), .ZN(new_n474));
  OR2_X1    g402(.A1(new_n330), .A2(new_n334), .ZN(new_n475));
  XOR2_X1   g403(.A(new_n470), .B(new_n471), .Z(new_n476));
  XOR2_X1   g404(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g405(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g406(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g407(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g408(.A(new_n480), .B1(new_n473), .B2(new_n479), .ZN(new_n481));
  INV_X1    g409(.A(new_n481), .ZN(new_n482));
  OAI221_X1 g410(.A(new_n469), .B1(new_n404), .B2(new_n473), .C1(new_n277), .C2(new_n482), .ZN(G3534));
  OAI21_X1  g411(.A(new_n216), .B1(new_n204), .B2(new_n265), .ZN(new_n484));
  INV_X1    g412(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g413(.A(new_n485), .B1(new_n215), .B2(new_n264), .ZN(new_n486));
  OR2_X1    g414(.A1(new_n364), .A2(new_n373), .ZN(new_n487));
  NAND2_X1  g415(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g416(.A(new_n281), .B1(new_n474), .B2(new_n478), .ZN(new_n489));
  INV_X1    g417(.A(new_n480), .ZN(new_n490));
  AOI21_X1  g418(.A(new_n489), .B1(new_n478), .B2(new_n490), .ZN(new_n491));
  OAI221_X1 g419(.A(new_n488), .B1(new_n486), .B2(new_n487), .C1(new_n283), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g420(.A1(new_n351), .A2(new_n486), .ZN(new_n493));
  OAI21_X1  g421(.A(new_n296), .B1(G15), .B2(G19), .ZN(new_n494));
  OAI211_X1 g422(.A(new_n143), .B(new_n494), .C1(new_n300), .C2(new_n342), .ZN(new_n495));
  AOI21_X1  g423(.A(new_n495), .B1(G21), .B2(new_n310), .ZN(new_n496));
  INV_X1    g424(.A(G17), .ZN(new_n497));
  AOI21_X1  g425(.A(G20), .B1(G16), .B2(new_n303), .ZN(new_n498));
  OAI221_X1 g426(.A(new_n496), .B1(new_n497), .B2(new_n311), .C1(new_n308), .C2(new_n498), .ZN(new_n499));
  AOI21_X1  g427(.A(new_n295), .B1(G11), .B2(new_n190), .ZN(new_n500));
  OAI21_X1  g428(.A(new_n429), .B1(G14), .B2(new_n302), .ZN(new_n501));
  NOR4_X1   g429(.A1(new_n142), .A2(new_n381), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  OAI21_X1  g430(.A(new_n502), .B1(G13), .B2(new_n311), .ZN(new_n503));
  OAI221_X1 g431(.A(new_n499), .B1(G5), .B2(G7), .C1(new_n427), .C2(new_n503), .ZN(new_n504));
  INV_X1    g432(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g433(.A(new_n284), .B1(new_n287), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g434(.A(new_n492), .B1(new_n493), .B2(new_n506), .ZN(G3535));
  OAI21_X1  g435(.A(new_n296), .B1(new_n78), .B2(G41), .ZN(new_n508));
  OAI21_X1  g436(.A(new_n508), .B1(G3), .B2(G12), .ZN(new_n509));
  AOI21_X1  g437(.A(new_n509), .B1(new_n89), .B2(new_n310), .ZN(new_n510));
  OAI221_X1 g438(.A(new_n510), .B1(G10), .B2(new_n300), .C1(new_n302), .C2(new_n391), .ZN(new_n511));
  OAI222_X1 g439(.A1(new_n347), .A2(new_n300), .B1(G7), .B2(new_n305), .C1(new_n458), .C2(new_n302), .ZN(new_n512));
  AOI21_X1  g440(.A(new_n295), .B1(new_n497), .B2(new_n199), .ZN(new_n513));
  NOR3_X1   g441(.A1(G4), .A2(new_n513), .A3(new_n428), .ZN(new_n514));
  OAI221_X1 g442(.A(new_n514), .B1(new_n345), .B2(new_n311), .C1(new_n224), .C2(new_n308), .ZN(new_n515));
  OAI22_X1  g443(.A1(new_n419), .A2(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g444(.A(new_n516), .ZN(new_n517));
  OAI221_X1 g445(.A(new_n284), .B1(new_n287), .B2(new_n517), .C1(new_n351), .C2(new_n470), .ZN(new_n518));
  INV_X1    g446(.A(new_n479), .ZN(new_n519));
  OAI221_X1 g447(.A(new_n518), .B1(new_n404), .B2(new_n477), .C1(new_n519), .C2(new_n489), .ZN(G3536));
  OR4_X1    g448(.A1(G3528), .A2(G3532), .A3(G3533), .A4(G3531), .ZN(new_n521));
  NOR2_X1   g449(.A1(G3534), .A2(G3535), .ZN(new_n522));
  INV_X1    g450(.A(new_n522), .ZN(new_n523));
  OR4_X1    g451(.A1(G3529), .A2(G3536), .A3(new_n521), .A4(new_n523), .ZN(G3537));
  NOR2_X1   g452(.A1(new_n263), .A2(new_n262), .ZN(new_n525));
  INV_X1    g453(.A(new_n525), .ZN(new_n526));
  OAI211_X1 g454(.A(G27), .B(G3537), .C1(new_n523), .C2(new_n526), .ZN(G3538));
  XNOR2_X1  g455(.A(G3529), .B(G3536), .ZN(new_n528));
  XOR2_X1   g456(.A(G3528), .B(G3532), .Z(new_n529));
  XNOR2_X1  g457(.A(G3531), .B(new_n529), .ZN(new_n530));
  AOI21_X1  g458(.A(new_n522), .B1(G3534), .B2(G3535), .ZN(new_n531));
  XNOR2_X1  g459(.A(G3533), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g460(.A(new_n530), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g461(.A(new_n528), .B(new_n533), .ZN(G3540));
  OAI22_X1  g462(.A1(new_n526), .A2(new_n531), .B1(G50), .B2(new_n525), .ZN(new_n535));
  XOR2_X1   g463(.A(G3540), .B(new_n535), .Z(G3539));
endmodule


