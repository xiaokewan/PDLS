// Benchmark "iscas85-original/c6288" written by ABC on Sat Nov 18 15:16:06 2023

module c6288  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32,
    G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32;
  output G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288;
  wire new_n65, new_n66, new_n68, new_n69, new_n70, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89, new_n90,
    new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97, new_n98,
    new_n99, new_n100, new_n101, new_n102, new_n104, new_n105, new_n106,
    new_n107, new_n108, new_n109, new_n110, new_n111, new_n112, new_n113,
    new_n114, new_n115, new_n116, new_n117, new_n118, new_n119, new_n120,
    new_n121, new_n122, new_n123, new_n124, new_n125, new_n126, new_n127,
    new_n128, new_n129, new_n130, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378, new_n379, new_n380, new_n381, new_n382, new_n383, new_n384,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1361, new_n1362, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1549, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1567, new_n1568, new_n1569, new_n1570,
    new_n1571, new_n1572, new_n1573, new_n1574, new_n1575, new_n1576,
    new_n1577, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1584, new_n1585, new_n1586, new_n1587, new_n1588,
    new_n1589, new_n1590, new_n1591, new_n1592, new_n1593, new_n1594,
    new_n1595, new_n1596, new_n1597, new_n1598, new_n1599, new_n1600,
    new_n1601, new_n1602, new_n1603, new_n1604, new_n1605, new_n1606,
    new_n1607, new_n1608, new_n1609, new_n1610, new_n1611, new_n1612,
    new_n1613, new_n1614, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1626, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1633, new_n1634, new_n1635, new_n1636, new_n1637,
    new_n1638, new_n1639, new_n1640, new_n1641, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1656, new_n1657, new_n1658, new_n1659, new_n1660, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1878, new_n1879, new_n1880, new_n1881, new_n1882,
    new_n1883, new_n1884, new_n1885, new_n1886, new_n1887, new_n1888,
    new_n1889, new_n1890, new_n1891, new_n1892, new_n1893, new_n1894,
    new_n1895, new_n1896, new_n1897, new_n1898, new_n1899, new_n1900,
    new_n1901, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924;
  INV_X1    g0000(.A(G1), .ZN(new_n65));
  INV_X1    g0001(.A(G17), .ZN(new_n66));
  NOR2_X1   g0002(.A1(new_n65), .A2(new_n66), .ZN(G6257));
  AOI22_X1  g0003(.A1(G2), .A2(G17), .B1(G1), .B2(G18), .ZN(new_n68));
  NAND3_X1  g0004(.A1(G2), .A2(G18), .A3(G6257), .ZN(new_n69));
  INV_X1    g0005(.A(new_n69), .ZN(new_n70));
  NOR2_X1   g0006(.A1(new_n68), .A2(new_n70), .ZN(G6258));
  INV_X1    g0007(.A(G19), .ZN(new_n72));
  NOR2_X1   g0008(.A1(new_n65), .A2(new_n72), .ZN(new_n73));
  AOI22_X1  g0009(.A1(G2), .A2(G18), .B1(G3), .B2(G17), .ZN(new_n74));
  INV_X1    g0010(.A(G2), .ZN(new_n75));
  INV_X1    g0011(.A(G3), .ZN(new_n76));
  INV_X1    g0012(.A(G18), .ZN(new_n77));
  NOR4_X1   g0013(.A1(new_n75), .A2(new_n66), .A3(new_n76), .A4(new_n77), .ZN(new_n78));
  OAI21_X1  g0014(.A(new_n69), .B1(new_n74), .B2(new_n78), .ZN(new_n79));
  OAI21_X1  g0015(.A(new_n79), .B1(new_n69), .B2(new_n78), .ZN(new_n80));
  NOR2_X1   g0016(.A1(new_n73), .A2(new_n80), .ZN(new_n81));
  AOI21_X1  g0017(.A(new_n81), .B1(new_n73), .B2(new_n80), .ZN(new_n82));
  INV_X1    g0018(.A(new_n82), .ZN(G6259));
  INV_X1    g0019(.A(G20), .ZN(new_n84));
  NOR2_X1   g0020(.A1(new_n65), .A2(new_n84), .ZN(new_n85));
  NOR2_X1   g0021(.A1(new_n75), .A2(new_n72), .ZN(new_n86));
  INV_X1    g0022(.A(new_n78), .ZN(new_n87));
  AOI22_X1  g0023(.A1(G3), .A2(G18), .B1(G4), .B2(G17), .ZN(new_n88));
  INV_X1    g0024(.A(G4), .ZN(new_n89));
  NOR4_X1   g0025(.A1(new_n76), .A2(new_n66), .A3(new_n89), .A4(new_n77), .ZN(new_n90));
  OAI21_X1  g0026(.A(new_n87), .B1(new_n88), .B2(new_n90), .ZN(new_n91));
  OAI21_X1  g0027(.A(new_n91), .B1(new_n87), .B2(new_n90), .ZN(new_n92));
  NOR2_X1   g0028(.A1(new_n86), .A2(new_n92), .ZN(new_n93));
  AOI21_X1  g0029(.A(new_n93), .B1(new_n86), .B2(new_n92), .ZN(new_n94));
  INV_X1    g0030(.A(new_n94), .ZN(new_n95));
  INV_X1    g0031(.A(new_n79), .ZN(new_n96));
  NOR2_X1   g0032(.A1(new_n96), .A2(new_n81), .ZN(new_n97));
  NOR2_X1   g0033(.A1(new_n95), .A2(new_n97), .ZN(new_n98));
  AOI21_X1  g0034(.A(new_n98), .B1(new_n95), .B2(new_n97), .ZN(new_n99));
  INV_X1    g0035(.A(new_n99), .ZN(new_n100));
  NOR2_X1   g0036(.A1(new_n85), .A2(new_n100), .ZN(new_n101));
  AOI21_X1  g0037(.A(new_n101), .B1(new_n85), .B2(new_n100), .ZN(new_n102));
  INV_X1    g0038(.A(new_n102), .ZN(G6260));
  INV_X1    g0039(.A(G21), .ZN(new_n104));
  NOR2_X1   g0040(.A1(new_n65), .A2(new_n104), .ZN(new_n105));
  NOR2_X1   g0041(.A1(new_n75), .A2(new_n84), .ZN(new_n106));
  NOR2_X1   g0042(.A1(new_n76), .A2(new_n72), .ZN(new_n107));
  INV_X1    g0043(.A(new_n90), .ZN(new_n108));
  AOI22_X1  g0044(.A1(G4), .A2(G18), .B1(G5), .B2(G17), .ZN(new_n109));
  INV_X1    g0045(.A(G5), .ZN(new_n110));
  NOR4_X1   g0046(.A1(new_n89), .A2(new_n66), .A3(new_n110), .A4(new_n77), .ZN(new_n111));
  OAI21_X1  g0047(.A(new_n108), .B1(new_n109), .B2(new_n111), .ZN(new_n112));
  OAI21_X1  g0048(.A(new_n112), .B1(new_n108), .B2(new_n111), .ZN(new_n113));
  NOR2_X1   g0049(.A1(new_n107), .A2(new_n113), .ZN(new_n114));
  AOI21_X1  g0050(.A(new_n114), .B1(new_n107), .B2(new_n113), .ZN(new_n115));
  INV_X1    g0051(.A(new_n115), .ZN(new_n116));
  INV_X1    g0052(.A(new_n91), .ZN(new_n117));
  NOR2_X1   g0053(.A1(new_n117), .A2(new_n93), .ZN(new_n118));
  NOR2_X1   g0054(.A1(new_n116), .A2(new_n118), .ZN(new_n119));
  AOI21_X1  g0055(.A(new_n119), .B1(new_n116), .B2(new_n118), .ZN(new_n120));
  INV_X1    g0056(.A(new_n120), .ZN(new_n121));
  NOR2_X1   g0057(.A1(new_n106), .A2(new_n121), .ZN(new_n122));
  AOI21_X1  g0058(.A(new_n122), .B1(new_n106), .B2(new_n121), .ZN(new_n123));
  INV_X1    g0059(.A(new_n123), .ZN(new_n124));
  NOR2_X1   g0060(.A1(new_n98), .A2(new_n101), .ZN(new_n125));
  NOR2_X1   g0061(.A1(new_n124), .A2(new_n125), .ZN(new_n126));
  AOI21_X1  g0062(.A(new_n126), .B1(new_n124), .B2(new_n125), .ZN(new_n127));
  INV_X1    g0063(.A(new_n127), .ZN(new_n128));
  NOR2_X1   g0064(.A1(new_n105), .A2(new_n128), .ZN(new_n129));
  AOI21_X1  g0065(.A(new_n129), .B1(new_n105), .B2(new_n128), .ZN(new_n130));
  INV_X1    g0066(.A(new_n130), .ZN(G6261));
  INV_X1    g0067(.A(G22), .ZN(new_n132));
  NOR2_X1   g0068(.A1(new_n65), .A2(new_n132), .ZN(new_n133));
  NOR2_X1   g0069(.A1(new_n75), .A2(new_n104), .ZN(new_n134));
  NOR2_X1   g0070(.A1(new_n76), .A2(new_n84), .ZN(new_n135));
  NOR2_X1   g0071(.A1(new_n89), .A2(new_n72), .ZN(new_n136));
  INV_X1    g0072(.A(new_n111), .ZN(new_n137));
  AOI22_X1  g0073(.A1(G5), .A2(G18), .B1(G6), .B2(G17), .ZN(new_n138));
  INV_X1    g0074(.A(G6), .ZN(new_n139));
  NOR4_X1   g0075(.A1(new_n110), .A2(new_n66), .A3(new_n139), .A4(new_n77), .ZN(new_n140));
  OAI21_X1  g0076(.A(new_n137), .B1(new_n138), .B2(new_n140), .ZN(new_n141));
  OAI21_X1  g0077(.A(new_n141), .B1(new_n137), .B2(new_n140), .ZN(new_n142));
  NOR2_X1   g0078(.A1(new_n136), .A2(new_n142), .ZN(new_n143));
  AOI21_X1  g0079(.A(new_n143), .B1(new_n136), .B2(new_n142), .ZN(new_n144));
  INV_X1    g0080(.A(new_n144), .ZN(new_n145));
  INV_X1    g0081(.A(new_n112), .ZN(new_n146));
  NOR2_X1   g0082(.A1(new_n146), .A2(new_n114), .ZN(new_n147));
  NOR2_X1   g0083(.A1(new_n145), .A2(new_n147), .ZN(new_n148));
  AOI21_X1  g0084(.A(new_n148), .B1(new_n145), .B2(new_n147), .ZN(new_n149));
  INV_X1    g0085(.A(new_n149), .ZN(new_n150));
  NOR2_X1   g0086(.A1(new_n135), .A2(new_n150), .ZN(new_n151));
  AOI21_X1  g0087(.A(new_n151), .B1(new_n135), .B2(new_n150), .ZN(new_n152));
  INV_X1    g0088(.A(new_n152), .ZN(new_n153));
  NOR2_X1   g0089(.A1(new_n119), .A2(new_n122), .ZN(new_n154));
  NOR2_X1   g0090(.A1(new_n153), .A2(new_n154), .ZN(new_n155));
  AOI21_X1  g0091(.A(new_n155), .B1(new_n153), .B2(new_n154), .ZN(new_n156));
  INV_X1    g0092(.A(new_n156), .ZN(new_n157));
  NOR2_X1   g0093(.A1(new_n134), .A2(new_n157), .ZN(new_n158));
  AOI21_X1  g0094(.A(new_n158), .B1(new_n134), .B2(new_n157), .ZN(new_n159));
  INV_X1    g0095(.A(new_n159), .ZN(new_n160));
  NOR2_X1   g0096(.A1(new_n126), .A2(new_n129), .ZN(new_n161));
  NOR2_X1   g0097(.A1(new_n160), .A2(new_n161), .ZN(new_n162));
  AOI21_X1  g0098(.A(new_n162), .B1(new_n160), .B2(new_n161), .ZN(new_n163));
  INV_X1    g0099(.A(new_n163), .ZN(new_n164));
  NOR2_X1   g0100(.A1(new_n133), .A2(new_n164), .ZN(new_n165));
  AOI21_X1  g0101(.A(new_n165), .B1(new_n133), .B2(new_n164), .ZN(new_n166));
  INV_X1    g0102(.A(new_n166), .ZN(G6262));
  INV_X1    g0103(.A(G23), .ZN(new_n168));
  NOR2_X1   g0104(.A1(new_n65), .A2(new_n168), .ZN(new_n169));
  NOR2_X1   g0105(.A1(new_n75), .A2(new_n132), .ZN(new_n170));
  NOR2_X1   g0106(.A1(new_n76), .A2(new_n104), .ZN(new_n171));
  NOR2_X1   g0107(.A1(new_n89), .A2(new_n84), .ZN(new_n172));
  NOR2_X1   g0108(.A1(new_n110), .A2(new_n72), .ZN(new_n173));
  INV_X1    g0109(.A(new_n140), .ZN(new_n174));
  AOI22_X1  g0110(.A1(G6), .A2(G18), .B1(G7), .B2(G17), .ZN(new_n175));
  INV_X1    g0111(.A(G7), .ZN(new_n176));
  NOR4_X1   g0112(.A1(new_n139), .A2(new_n66), .A3(new_n176), .A4(new_n77), .ZN(new_n177));
  OAI21_X1  g0113(.A(new_n174), .B1(new_n175), .B2(new_n177), .ZN(new_n178));
  OAI21_X1  g0114(.A(new_n178), .B1(new_n174), .B2(new_n177), .ZN(new_n179));
  NOR2_X1   g0115(.A1(new_n173), .A2(new_n179), .ZN(new_n180));
  AOI21_X1  g0116(.A(new_n180), .B1(new_n173), .B2(new_n179), .ZN(new_n181));
  INV_X1    g0117(.A(new_n181), .ZN(new_n182));
  INV_X1    g0118(.A(new_n141), .ZN(new_n183));
  NOR2_X1   g0119(.A1(new_n183), .A2(new_n143), .ZN(new_n184));
  NOR2_X1   g0120(.A1(new_n182), .A2(new_n184), .ZN(new_n185));
  AOI21_X1  g0121(.A(new_n185), .B1(new_n182), .B2(new_n184), .ZN(new_n186));
  INV_X1    g0122(.A(new_n186), .ZN(new_n187));
  NOR2_X1   g0123(.A1(new_n172), .A2(new_n187), .ZN(new_n188));
  AOI21_X1  g0124(.A(new_n188), .B1(new_n172), .B2(new_n187), .ZN(new_n189));
  INV_X1    g0125(.A(new_n189), .ZN(new_n190));
  NOR2_X1   g0126(.A1(new_n148), .A2(new_n151), .ZN(new_n191));
  NOR2_X1   g0127(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  AOI21_X1  g0128(.A(new_n192), .B1(new_n190), .B2(new_n191), .ZN(new_n193));
  INV_X1    g0129(.A(new_n193), .ZN(new_n194));
  NOR2_X1   g0130(.A1(new_n171), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g0131(.A(new_n195), .B1(new_n171), .B2(new_n194), .ZN(new_n196));
  INV_X1    g0132(.A(new_n196), .ZN(new_n197));
  NOR2_X1   g0133(.A1(new_n155), .A2(new_n158), .ZN(new_n198));
  NOR2_X1   g0134(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g0135(.A(new_n199), .B1(new_n197), .B2(new_n198), .ZN(new_n200));
  INV_X1    g0136(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g0137(.A1(new_n170), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g0138(.A(new_n202), .B1(new_n170), .B2(new_n201), .ZN(new_n203));
  INV_X1    g0139(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g0140(.A1(new_n162), .A2(new_n165), .ZN(new_n205));
  NOR2_X1   g0141(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g0142(.A(new_n206), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  INV_X1    g0143(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0144(.A1(new_n169), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g0145(.A(new_n209), .B1(new_n169), .B2(new_n208), .ZN(new_n210));
  INV_X1    g0146(.A(new_n210), .ZN(G6263));
  INV_X1    g0147(.A(G24), .ZN(new_n212));
  NOR2_X1   g0148(.A1(new_n65), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g0149(.A1(new_n75), .A2(new_n168), .ZN(new_n214));
  NOR2_X1   g0150(.A1(new_n76), .A2(new_n132), .ZN(new_n215));
  NOR2_X1   g0151(.A1(new_n89), .A2(new_n104), .ZN(new_n216));
  NOR2_X1   g0152(.A1(new_n110), .A2(new_n84), .ZN(new_n217));
  NOR2_X1   g0153(.A1(new_n139), .A2(new_n72), .ZN(new_n218));
  INV_X1    g0154(.A(new_n177), .ZN(new_n219));
  AOI22_X1  g0155(.A1(G7), .A2(G18), .B1(G8), .B2(G17), .ZN(new_n220));
  INV_X1    g0156(.A(G8), .ZN(new_n221));
  NOR4_X1   g0157(.A1(new_n176), .A2(new_n66), .A3(new_n221), .A4(new_n77), .ZN(new_n222));
  OAI21_X1  g0158(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g0159(.A(new_n223), .B1(new_n219), .B2(new_n222), .ZN(new_n224));
  NOR2_X1   g0160(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g0161(.A(new_n225), .B1(new_n218), .B2(new_n224), .ZN(new_n226));
  INV_X1    g0162(.A(new_n226), .ZN(new_n227));
  INV_X1    g0163(.A(new_n178), .ZN(new_n228));
  NOR2_X1   g0164(.A1(new_n228), .A2(new_n180), .ZN(new_n229));
  NOR2_X1   g0165(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g0166(.A(new_n230), .B1(new_n227), .B2(new_n229), .ZN(new_n231));
  INV_X1    g0167(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g0168(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g0169(.A(new_n233), .B1(new_n217), .B2(new_n232), .ZN(new_n234));
  INV_X1    g0170(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g0171(.A1(new_n185), .A2(new_n188), .ZN(new_n236));
  NOR2_X1   g0172(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g0173(.A(new_n237), .B1(new_n235), .B2(new_n236), .ZN(new_n238));
  INV_X1    g0174(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g0175(.A1(new_n216), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g0176(.A(new_n240), .B1(new_n216), .B2(new_n239), .ZN(new_n241));
  INV_X1    g0177(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g0178(.A1(new_n192), .A2(new_n195), .ZN(new_n243));
  NOR2_X1   g0179(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g0180(.A(new_n244), .B1(new_n242), .B2(new_n243), .ZN(new_n245));
  INV_X1    g0181(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g0182(.A1(new_n215), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g0183(.A(new_n247), .B1(new_n215), .B2(new_n246), .ZN(new_n248));
  INV_X1    g0184(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g0185(.A1(new_n199), .A2(new_n202), .ZN(new_n250));
  NOR2_X1   g0186(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g0187(.A(new_n251), .B1(new_n249), .B2(new_n250), .ZN(new_n252));
  INV_X1    g0188(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0189(.A1(new_n214), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0190(.A(new_n254), .B1(new_n214), .B2(new_n253), .ZN(new_n255));
  INV_X1    g0191(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0192(.A1(new_n206), .A2(new_n209), .ZN(new_n257));
  NOR2_X1   g0193(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0194(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n259));
  INV_X1    g0195(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0196(.A1(new_n213), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0197(.A(new_n261), .B1(new_n213), .B2(new_n260), .ZN(new_n262));
  INV_X1    g0198(.A(new_n262), .ZN(G6264));
  INV_X1    g0199(.A(G25), .ZN(new_n264));
  NOR2_X1   g0200(.A1(new_n65), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0201(.A1(new_n75), .A2(new_n212), .ZN(new_n266));
  NOR2_X1   g0202(.A1(new_n76), .A2(new_n168), .ZN(new_n267));
  NOR2_X1   g0203(.A1(new_n89), .A2(new_n132), .ZN(new_n268));
  NOR2_X1   g0204(.A1(new_n110), .A2(new_n104), .ZN(new_n269));
  NOR2_X1   g0205(.A1(new_n139), .A2(new_n84), .ZN(new_n270));
  NOR2_X1   g0206(.A1(new_n176), .A2(new_n72), .ZN(new_n271));
  INV_X1    g0207(.A(new_n222), .ZN(new_n272));
  AOI22_X1  g0208(.A1(G8), .A2(G18), .B1(G9), .B2(G17), .ZN(new_n273));
  INV_X1    g0209(.A(G9), .ZN(new_n274));
  NOR4_X1   g0210(.A1(new_n221), .A2(new_n66), .A3(new_n274), .A4(new_n77), .ZN(new_n275));
  OAI21_X1  g0211(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0212(.A(new_n276), .B1(new_n272), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g0213(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0214(.A(new_n278), .B1(new_n271), .B2(new_n277), .ZN(new_n279));
  INV_X1    g0215(.A(new_n279), .ZN(new_n280));
  INV_X1    g0216(.A(new_n223), .ZN(new_n281));
  NOR2_X1   g0217(.A1(new_n281), .A2(new_n225), .ZN(new_n282));
  NOR2_X1   g0218(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0219(.A(new_n283), .B1(new_n280), .B2(new_n282), .ZN(new_n284));
  INV_X1    g0220(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0221(.A1(new_n270), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0222(.A(new_n286), .B1(new_n270), .B2(new_n285), .ZN(new_n287));
  INV_X1    g0223(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0224(.A1(new_n230), .A2(new_n233), .ZN(new_n289));
  NOR2_X1   g0225(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0226(.A(new_n290), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  INV_X1    g0227(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0228(.A1(new_n269), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0229(.A(new_n293), .B1(new_n269), .B2(new_n292), .ZN(new_n294));
  INV_X1    g0230(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0231(.A1(new_n237), .A2(new_n240), .ZN(new_n296));
  NOR2_X1   g0232(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0233(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  INV_X1    g0234(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0235(.A1(new_n268), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0236(.A(new_n300), .B1(new_n268), .B2(new_n299), .ZN(new_n301));
  INV_X1    g0237(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0238(.A1(new_n244), .A2(new_n247), .ZN(new_n303));
  NOR2_X1   g0239(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0240(.A(new_n304), .B1(new_n302), .B2(new_n303), .ZN(new_n305));
  INV_X1    g0241(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0242(.A1(new_n267), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0243(.A(new_n307), .B1(new_n267), .B2(new_n306), .ZN(new_n308));
  INV_X1    g0244(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g0245(.A1(new_n251), .A2(new_n254), .ZN(new_n310));
  NOR2_X1   g0246(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0247(.A(new_n311), .B1(new_n309), .B2(new_n310), .ZN(new_n312));
  INV_X1    g0248(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g0249(.A1(new_n266), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0250(.A(new_n314), .B1(new_n266), .B2(new_n313), .ZN(new_n315));
  INV_X1    g0251(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0252(.A1(new_n258), .A2(new_n261), .ZN(new_n317));
  NOR2_X1   g0253(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0254(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  INV_X1    g0255(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g0256(.A1(new_n265), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0257(.A(new_n321), .B1(new_n265), .B2(new_n320), .ZN(new_n322));
  INV_X1    g0258(.A(new_n322), .ZN(G6265));
  INV_X1    g0259(.A(G26), .ZN(new_n324));
  NOR2_X1   g0260(.A1(new_n65), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0261(.A1(new_n75), .A2(new_n264), .ZN(new_n326));
  NOR2_X1   g0262(.A1(new_n76), .A2(new_n212), .ZN(new_n327));
  NOR2_X1   g0263(.A1(new_n89), .A2(new_n168), .ZN(new_n328));
  NOR2_X1   g0264(.A1(new_n110), .A2(new_n132), .ZN(new_n329));
  NOR2_X1   g0265(.A1(new_n139), .A2(new_n104), .ZN(new_n330));
  NOR2_X1   g0266(.A1(new_n176), .A2(new_n84), .ZN(new_n331));
  NOR2_X1   g0267(.A1(new_n221), .A2(new_n72), .ZN(new_n332));
  INV_X1    g0268(.A(new_n275), .ZN(new_n333));
  AOI22_X1  g0269(.A1(G9), .A2(G18), .B1(G10), .B2(G17), .ZN(new_n334));
  INV_X1    g0270(.A(G10), .ZN(new_n335));
  NOR4_X1   g0271(.A1(new_n274), .A2(new_n66), .A3(new_n335), .A4(new_n77), .ZN(new_n336));
  OAI21_X1  g0272(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0273(.A(new_n337), .B1(new_n333), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0274(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0275(.A(new_n339), .B1(new_n332), .B2(new_n338), .ZN(new_n340));
  INV_X1    g0276(.A(new_n340), .ZN(new_n341));
  INV_X1    g0277(.A(new_n276), .ZN(new_n342));
  NOR2_X1   g0278(.A1(new_n342), .A2(new_n278), .ZN(new_n343));
  NOR2_X1   g0279(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0280(.A(new_n344), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  INV_X1    g0281(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g0282(.A1(new_n331), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0283(.A(new_n347), .B1(new_n331), .B2(new_n346), .ZN(new_n348));
  INV_X1    g0284(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g0285(.A1(new_n283), .A2(new_n286), .ZN(new_n350));
  NOR2_X1   g0286(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0287(.A(new_n351), .B1(new_n349), .B2(new_n350), .ZN(new_n352));
  INV_X1    g0288(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g0289(.A1(new_n330), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0290(.A(new_n354), .B1(new_n330), .B2(new_n353), .ZN(new_n355));
  INV_X1    g0291(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0292(.A1(new_n290), .A2(new_n293), .ZN(new_n357));
  NOR2_X1   g0293(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0294(.A(new_n358), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  INV_X1    g0295(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0296(.A1(new_n329), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0297(.A(new_n361), .B1(new_n329), .B2(new_n360), .ZN(new_n362));
  INV_X1    g0298(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0299(.A1(new_n297), .A2(new_n300), .ZN(new_n364));
  NOR2_X1   g0300(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0301(.A(new_n365), .B1(new_n363), .B2(new_n364), .ZN(new_n366));
  INV_X1    g0302(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g0303(.A1(new_n328), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0304(.A(new_n368), .B1(new_n328), .B2(new_n367), .ZN(new_n369));
  INV_X1    g0305(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g0306(.A1(new_n304), .A2(new_n307), .ZN(new_n371));
  NOR2_X1   g0307(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0308(.A(new_n372), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  INV_X1    g0309(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g0310(.A1(new_n327), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0311(.A(new_n375), .B1(new_n327), .B2(new_n374), .ZN(new_n376));
  INV_X1    g0312(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0313(.A1(new_n311), .A2(new_n314), .ZN(new_n378));
  NOR2_X1   g0314(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0315(.A(new_n379), .B1(new_n377), .B2(new_n378), .ZN(new_n380));
  INV_X1    g0316(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g0317(.A1(new_n326), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0318(.A(new_n382), .B1(new_n326), .B2(new_n381), .ZN(new_n383));
  INV_X1    g0319(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0320(.A1(new_n318), .A2(new_n321), .ZN(new_n385));
  NOR2_X1   g0321(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0322(.A(new_n386), .B1(new_n384), .B2(new_n385), .ZN(new_n387));
  INV_X1    g0323(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g0324(.A1(new_n325), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0325(.A(new_n389), .B1(new_n325), .B2(new_n388), .ZN(new_n390));
  INV_X1    g0326(.A(new_n390), .ZN(G6266));
  INV_X1    g0327(.A(G27), .ZN(new_n392));
  NOR2_X1   g0328(.A1(new_n65), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0329(.A1(new_n75), .A2(new_n324), .ZN(new_n394));
  NOR2_X1   g0330(.A1(new_n76), .A2(new_n264), .ZN(new_n395));
  NOR2_X1   g0331(.A1(new_n89), .A2(new_n212), .ZN(new_n396));
  NOR2_X1   g0332(.A1(new_n110), .A2(new_n168), .ZN(new_n397));
  NOR2_X1   g0333(.A1(new_n139), .A2(new_n132), .ZN(new_n398));
  NOR2_X1   g0334(.A1(new_n176), .A2(new_n104), .ZN(new_n399));
  NOR2_X1   g0335(.A1(new_n221), .A2(new_n84), .ZN(new_n400));
  NOR2_X1   g0336(.A1(new_n274), .A2(new_n72), .ZN(new_n401));
  INV_X1    g0337(.A(new_n336), .ZN(new_n402));
  AOI22_X1  g0338(.A1(G10), .A2(G18), .B1(G11), .B2(G17), .ZN(new_n403));
  INV_X1    g0339(.A(G11), .ZN(new_n404));
  NOR4_X1   g0340(.A1(new_n335), .A2(new_n66), .A3(new_n404), .A4(new_n77), .ZN(new_n405));
  OAI21_X1  g0341(.A(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0342(.A(new_n406), .B1(new_n402), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g0343(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0344(.A(new_n408), .B1(new_n401), .B2(new_n407), .ZN(new_n409));
  INV_X1    g0345(.A(new_n409), .ZN(new_n410));
  INV_X1    g0346(.A(new_n337), .ZN(new_n411));
  NOR2_X1   g0347(.A1(new_n411), .A2(new_n339), .ZN(new_n412));
  NOR2_X1   g0348(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0349(.A(new_n413), .B1(new_n410), .B2(new_n412), .ZN(new_n414));
  INV_X1    g0350(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g0351(.A1(new_n400), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0352(.A(new_n416), .B1(new_n400), .B2(new_n415), .ZN(new_n417));
  INV_X1    g0353(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g0354(.A1(new_n344), .A2(new_n347), .ZN(new_n419));
  NOR2_X1   g0355(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0356(.A(new_n420), .B1(new_n418), .B2(new_n419), .ZN(new_n421));
  INV_X1    g0357(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0358(.A1(new_n399), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0359(.A(new_n423), .B1(new_n399), .B2(new_n422), .ZN(new_n424));
  INV_X1    g0360(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g0361(.A1(new_n351), .A2(new_n354), .ZN(new_n426));
  NOR2_X1   g0362(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0363(.A(new_n427), .B1(new_n425), .B2(new_n426), .ZN(new_n428));
  INV_X1    g0364(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g0365(.A1(new_n398), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0366(.A(new_n430), .B1(new_n398), .B2(new_n429), .ZN(new_n431));
  INV_X1    g0367(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g0368(.A1(new_n358), .A2(new_n361), .ZN(new_n433));
  NOR2_X1   g0369(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0370(.A(new_n434), .B1(new_n432), .B2(new_n433), .ZN(new_n435));
  INV_X1    g0371(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0372(.A1(new_n397), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0373(.A(new_n437), .B1(new_n397), .B2(new_n436), .ZN(new_n438));
  INV_X1    g0374(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g0375(.A1(new_n365), .A2(new_n368), .ZN(new_n440));
  NOR2_X1   g0376(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0377(.A(new_n441), .B1(new_n439), .B2(new_n440), .ZN(new_n442));
  INV_X1    g0378(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g0379(.A1(new_n396), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0380(.A(new_n444), .B1(new_n396), .B2(new_n443), .ZN(new_n445));
  INV_X1    g0381(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g0382(.A1(new_n372), .A2(new_n375), .ZN(new_n447));
  NOR2_X1   g0383(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0384(.A(new_n448), .B1(new_n446), .B2(new_n447), .ZN(new_n449));
  INV_X1    g0385(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g0386(.A1(new_n395), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0387(.A(new_n451), .B1(new_n395), .B2(new_n450), .ZN(new_n452));
  INV_X1    g0388(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g0389(.A1(new_n379), .A2(new_n382), .ZN(new_n454));
  NOR2_X1   g0390(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0391(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n456));
  INV_X1    g0392(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0393(.A1(new_n394), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0394(.A(new_n458), .B1(new_n394), .B2(new_n457), .ZN(new_n459));
  INV_X1    g0395(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0396(.A1(new_n386), .A2(new_n389), .ZN(new_n461));
  NOR2_X1   g0397(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0398(.A(new_n462), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  INV_X1    g0399(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g0400(.A1(new_n393), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0401(.A(new_n465), .B1(new_n393), .B2(new_n464), .ZN(new_n466));
  INV_X1    g0402(.A(new_n466), .ZN(G6267));
  INV_X1    g0403(.A(G28), .ZN(new_n468));
  NOR2_X1   g0404(.A1(new_n65), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0405(.A1(new_n75), .A2(new_n392), .ZN(new_n470));
  NOR2_X1   g0406(.A1(new_n76), .A2(new_n324), .ZN(new_n471));
  NOR2_X1   g0407(.A1(new_n89), .A2(new_n264), .ZN(new_n472));
  NOR2_X1   g0408(.A1(new_n110), .A2(new_n212), .ZN(new_n473));
  NOR2_X1   g0409(.A1(new_n139), .A2(new_n168), .ZN(new_n474));
  NOR2_X1   g0410(.A1(new_n176), .A2(new_n132), .ZN(new_n475));
  NOR2_X1   g0411(.A1(new_n221), .A2(new_n104), .ZN(new_n476));
  NOR2_X1   g0412(.A1(new_n274), .A2(new_n84), .ZN(new_n477));
  NOR2_X1   g0413(.A1(new_n335), .A2(new_n72), .ZN(new_n478));
  INV_X1    g0414(.A(new_n405), .ZN(new_n479));
  AOI22_X1  g0415(.A1(G11), .A2(G18), .B1(G12), .B2(G17), .ZN(new_n480));
  INV_X1    g0416(.A(G12), .ZN(new_n481));
  NOR4_X1   g0417(.A1(new_n404), .A2(new_n66), .A3(new_n481), .A4(new_n77), .ZN(new_n482));
  OAI21_X1  g0418(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0419(.A(new_n483), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g0420(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0421(.A(new_n485), .B1(new_n478), .B2(new_n484), .ZN(new_n486));
  INV_X1    g0422(.A(new_n486), .ZN(new_n487));
  INV_X1    g0423(.A(new_n406), .ZN(new_n488));
  NOR2_X1   g0424(.A1(new_n488), .A2(new_n408), .ZN(new_n489));
  NOR2_X1   g0425(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0426(.A(new_n490), .B1(new_n487), .B2(new_n489), .ZN(new_n491));
  INV_X1    g0427(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g0428(.A1(new_n477), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0429(.A(new_n493), .B1(new_n477), .B2(new_n492), .ZN(new_n494));
  INV_X1    g0430(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0431(.A1(new_n413), .A2(new_n416), .ZN(new_n496));
  NOR2_X1   g0432(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0433(.A(new_n497), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  INV_X1    g0434(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g0435(.A1(new_n476), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0436(.A(new_n500), .B1(new_n476), .B2(new_n499), .ZN(new_n501));
  INV_X1    g0437(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0438(.A1(new_n420), .A2(new_n423), .ZN(new_n503));
  NOR2_X1   g0439(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0440(.A(new_n504), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  INV_X1    g0441(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0442(.A1(new_n475), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0443(.A(new_n507), .B1(new_n475), .B2(new_n506), .ZN(new_n508));
  INV_X1    g0444(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0445(.A1(new_n427), .A2(new_n430), .ZN(new_n510));
  NOR2_X1   g0446(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0447(.A(new_n511), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  INV_X1    g0448(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0449(.A1(new_n474), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0450(.A(new_n514), .B1(new_n474), .B2(new_n513), .ZN(new_n515));
  INV_X1    g0451(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g0452(.A1(new_n434), .A2(new_n437), .ZN(new_n517));
  NOR2_X1   g0453(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0454(.A(new_n518), .B1(new_n516), .B2(new_n517), .ZN(new_n519));
  INV_X1    g0455(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g0456(.A1(new_n473), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0457(.A(new_n521), .B1(new_n473), .B2(new_n520), .ZN(new_n522));
  INV_X1    g0458(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g0459(.A1(new_n441), .A2(new_n444), .ZN(new_n524));
  NOR2_X1   g0460(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0461(.A(new_n525), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  INV_X1    g0462(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g0463(.A1(new_n472), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0464(.A(new_n528), .B1(new_n472), .B2(new_n527), .ZN(new_n529));
  INV_X1    g0465(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g0466(.A1(new_n448), .A2(new_n451), .ZN(new_n531));
  NOR2_X1   g0467(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0468(.A(new_n532), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  INV_X1    g0469(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g0470(.A1(new_n471), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0471(.A(new_n535), .B1(new_n471), .B2(new_n534), .ZN(new_n536));
  INV_X1    g0472(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0473(.A1(new_n455), .A2(new_n458), .ZN(new_n538));
  NOR2_X1   g0474(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0475(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n540));
  INV_X1    g0476(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g0477(.A1(new_n470), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0478(.A(new_n542), .B1(new_n470), .B2(new_n541), .ZN(new_n543));
  INV_X1    g0479(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0480(.A1(new_n462), .A2(new_n465), .ZN(new_n545));
  NOR2_X1   g0481(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0482(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  INV_X1    g0483(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g0484(.A1(new_n469), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0485(.A(new_n549), .B1(new_n469), .B2(new_n548), .ZN(new_n550));
  INV_X1    g0486(.A(new_n550), .ZN(G6268));
  INV_X1    g0487(.A(G29), .ZN(new_n552));
  NOR2_X1   g0488(.A1(new_n65), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0489(.A1(new_n75), .A2(new_n468), .ZN(new_n554));
  NOR2_X1   g0490(.A1(new_n76), .A2(new_n392), .ZN(new_n555));
  NOR2_X1   g0491(.A1(new_n89), .A2(new_n324), .ZN(new_n556));
  NOR2_X1   g0492(.A1(new_n110), .A2(new_n264), .ZN(new_n557));
  NOR2_X1   g0493(.A1(new_n139), .A2(new_n212), .ZN(new_n558));
  NOR2_X1   g0494(.A1(new_n176), .A2(new_n168), .ZN(new_n559));
  NOR2_X1   g0495(.A1(new_n221), .A2(new_n132), .ZN(new_n560));
  NOR2_X1   g0496(.A1(new_n274), .A2(new_n104), .ZN(new_n561));
  NOR2_X1   g0497(.A1(new_n335), .A2(new_n84), .ZN(new_n562));
  NOR2_X1   g0498(.A1(new_n404), .A2(new_n72), .ZN(new_n563));
  INV_X1    g0499(.A(new_n482), .ZN(new_n564));
  AOI22_X1  g0500(.A1(G12), .A2(G18), .B1(G13), .B2(G17), .ZN(new_n565));
  INV_X1    g0501(.A(G13), .ZN(new_n566));
  NOR4_X1   g0502(.A1(new_n481), .A2(new_n66), .A3(new_n566), .A4(new_n77), .ZN(new_n567));
  OAI21_X1  g0503(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0504(.A(new_n568), .B1(new_n564), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g0505(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0506(.A(new_n570), .B1(new_n563), .B2(new_n569), .ZN(new_n571));
  INV_X1    g0507(.A(new_n571), .ZN(new_n572));
  INV_X1    g0508(.A(new_n483), .ZN(new_n573));
  NOR2_X1   g0509(.A1(new_n573), .A2(new_n485), .ZN(new_n574));
  NOR2_X1   g0510(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0511(.A(new_n575), .B1(new_n572), .B2(new_n574), .ZN(new_n576));
  INV_X1    g0512(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g0513(.A1(new_n562), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0514(.A(new_n578), .B1(new_n562), .B2(new_n577), .ZN(new_n579));
  INV_X1    g0515(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g0516(.A1(new_n490), .A2(new_n493), .ZN(new_n581));
  NOR2_X1   g0517(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0518(.A(new_n582), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  INV_X1    g0519(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g0520(.A1(new_n561), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0521(.A(new_n585), .B1(new_n561), .B2(new_n584), .ZN(new_n586));
  INV_X1    g0522(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g0523(.A1(new_n497), .A2(new_n500), .ZN(new_n588));
  NOR2_X1   g0524(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0525(.A(new_n589), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  INV_X1    g0526(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g0527(.A1(new_n560), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0528(.A(new_n592), .B1(new_n560), .B2(new_n591), .ZN(new_n593));
  INV_X1    g0529(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g0530(.A1(new_n504), .A2(new_n507), .ZN(new_n595));
  NOR2_X1   g0531(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0532(.A(new_n596), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  INV_X1    g0533(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g0534(.A1(new_n559), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0535(.A(new_n599), .B1(new_n559), .B2(new_n598), .ZN(new_n600));
  INV_X1    g0536(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g0537(.A1(new_n511), .A2(new_n514), .ZN(new_n602));
  NOR2_X1   g0538(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0539(.A(new_n603), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  INV_X1    g0540(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g0541(.A1(new_n558), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0542(.A(new_n606), .B1(new_n558), .B2(new_n605), .ZN(new_n607));
  INV_X1    g0543(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g0544(.A1(new_n518), .A2(new_n521), .ZN(new_n609));
  NOR2_X1   g0545(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0546(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  INV_X1    g0547(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g0548(.A1(new_n557), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0549(.A(new_n613), .B1(new_n557), .B2(new_n612), .ZN(new_n614));
  INV_X1    g0550(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g0551(.A1(new_n525), .A2(new_n528), .ZN(new_n616));
  NOR2_X1   g0552(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0553(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  INV_X1    g0554(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g0555(.A1(new_n556), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0556(.A(new_n620), .B1(new_n556), .B2(new_n619), .ZN(new_n621));
  INV_X1    g0557(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0558(.A1(new_n532), .A2(new_n535), .ZN(new_n623));
  NOR2_X1   g0559(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0560(.A(new_n624), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  INV_X1    g0561(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0562(.A1(new_n555), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0563(.A(new_n627), .B1(new_n555), .B2(new_n626), .ZN(new_n628));
  INV_X1    g0564(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g0565(.A1(new_n539), .A2(new_n542), .ZN(new_n630));
  NOR2_X1   g0566(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0567(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  INV_X1    g0568(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g0569(.A1(new_n554), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0570(.A(new_n634), .B1(new_n554), .B2(new_n633), .ZN(new_n635));
  INV_X1    g0571(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0572(.A1(new_n546), .A2(new_n549), .ZN(new_n637));
  NOR2_X1   g0573(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0574(.A(new_n638), .B1(new_n636), .B2(new_n637), .ZN(new_n639));
  INV_X1    g0575(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0576(.A1(new_n553), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0577(.A(new_n641), .B1(new_n553), .B2(new_n640), .ZN(new_n642));
  INV_X1    g0578(.A(new_n642), .ZN(G6269));
  INV_X1    g0579(.A(G30), .ZN(new_n644));
  NOR2_X1   g0580(.A1(new_n65), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0581(.A1(new_n75), .A2(new_n552), .ZN(new_n646));
  NOR2_X1   g0582(.A1(new_n76), .A2(new_n468), .ZN(new_n647));
  NOR2_X1   g0583(.A1(new_n89), .A2(new_n392), .ZN(new_n648));
  NOR2_X1   g0584(.A1(new_n110), .A2(new_n324), .ZN(new_n649));
  NOR2_X1   g0585(.A1(new_n139), .A2(new_n264), .ZN(new_n650));
  NOR2_X1   g0586(.A1(new_n176), .A2(new_n212), .ZN(new_n651));
  NOR2_X1   g0587(.A1(new_n221), .A2(new_n168), .ZN(new_n652));
  NOR2_X1   g0588(.A1(new_n274), .A2(new_n132), .ZN(new_n653));
  NOR2_X1   g0589(.A1(new_n335), .A2(new_n104), .ZN(new_n654));
  NOR2_X1   g0590(.A1(new_n404), .A2(new_n84), .ZN(new_n655));
  NOR2_X1   g0591(.A1(new_n481), .A2(new_n72), .ZN(new_n656));
  INV_X1    g0592(.A(new_n567), .ZN(new_n657));
  AOI22_X1  g0593(.A1(G13), .A2(G18), .B1(G14), .B2(G17), .ZN(new_n658));
  INV_X1    g0594(.A(G14), .ZN(new_n659));
  NOR4_X1   g0595(.A1(new_n566), .A2(new_n66), .A3(new_n659), .A4(new_n77), .ZN(new_n660));
  OAI21_X1  g0596(.A(new_n657), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0597(.A(new_n661), .B1(new_n657), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0598(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0599(.A(new_n663), .B1(new_n656), .B2(new_n662), .ZN(new_n664));
  INV_X1    g0600(.A(new_n664), .ZN(new_n665));
  INV_X1    g0601(.A(new_n568), .ZN(new_n666));
  NOR2_X1   g0602(.A1(new_n666), .A2(new_n570), .ZN(new_n667));
  NOR2_X1   g0603(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0604(.A(new_n668), .B1(new_n665), .B2(new_n667), .ZN(new_n669));
  INV_X1    g0605(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0606(.A1(new_n655), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0607(.A(new_n671), .B1(new_n655), .B2(new_n670), .ZN(new_n672));
  INV_X1    g0608(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0609(.A1(new_n575), .A2(new_n578), .ZN(new_n674));
  NOR2_X1   g0610(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0611(.A(new_n675), .B1(new_n673), .B2(new_n674), .ZN(new_n676));
  INV_X1    g0612(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0613(.A1(new_n654), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0614(.A(new_n678), .B1(new_n654), .B2(new_n677), .ZN(new_n679));
  INV_X1    g0615(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0616(.A1(new_n582), .A2(new_n585), .ZN(new_n681));
  NOR2_X1   g0617(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0618(.A(new_n682), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  INV_X1    g0619(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0620(.A1(new_n653), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0621(.A(new_n685), .B1(new_n653), .B2(new_n684), .ZN(new_n686));
  INV_X1    g0622(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0623(.A1(new_n589), .A2(new_n592), .ZN(new_n688));
  NOR2_X1   g0624(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0625(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  INV_X1    g0626(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0627(.A1(new_n652), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0628(.A(new_n692), .B1(new_n652), .B2(new_n691), .ZN(new_n693));
  INV_X1    g0629(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0630(.A1(new_n596), .A2(new_n599), .ZN(new_n695));
  NOR2_X1   g0631(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0632(.A(new_n696), .B1(new_n694), .B2(new_n695), .ZN(new_n697));
  INV_X1    g0633(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0634(.A1(new_n651), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0635(.A(new_n699), .B1(new_n651), .B2(new_n698), .ZN(new_n700));
  INV_X1    g0636(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0637(.A1(new_n603), .A2(new_n606), .ZN(new_n702));
  NOR2_X1   g0638(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0639(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  INV_X1    g0640(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0641(.A1(new_n650), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0642(.A(new_n706), .B1(new_n650), .B2(new_n705), .ZN(new_n707));
  INV_X1    g0643(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0644(.A1(new_n610), .A2(new_n613), .ZN(new_n709));
  NOR2_X1   g0645(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0646(.A(new_n710), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  INV_X1    g0647(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0648(.A1(new_n649), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0649(.A(new_n713), .B1(new_n649), .B2(new_n712), .ZN(new_n714));
  INV_X1    g0650(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0651(.A1(new_n617), .A2(new_n620), .ZN(new_n716));
  NOR2_X1   g0652(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0653(.A(new_n717), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  INV_X1    g0654(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0655(.A1(new_n648), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0656(.A(new_n720), .B1(new_n648), .B2(new_n719), .ZN(new_n721));
  INV_X1    g0657(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0658(.A1(new_n624), .A2(new_n627), .ZN(new_n723));
  NOR2_X1   g0659(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0660(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  INV_X1    g0661(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0662(.A1(new_n647), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0663(.A(new_n727), .B1(new_n647), .B2(new_n726), .ZN(new_n728));
  INV_X1    g0664(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0665(.A1(new_n631), .A2(new_n634), .ZN(new_n730));
  NOR2_X1   g0666(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0667(.A(new_n731), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  INV_X1    g0668(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0669(.A1(new_n646), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0670(.A(new_n734), .B1(new_n646), .B2(new_n733), .ZN(new_n735));
  INV_X1    g0671(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0672(.A1(new_n638), .A2(new_n641), .ZN(new_n737));
  NOR2_X1   g0673(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0674(.A(new_n738), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  INV_X1    g0675(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0676(.A1(new_n645), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0677(.A(new_n741), .B1(new_n645), .B2(new_n740), .ZN(new_n742));
  INV_X1    g0678(.A(new_n742), .ZN(G6270));
  INV_X1    g0679(.A(G31), .ZN(new_n744));
  NOR2_X1   g0680(.A1(new_n65), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0681(.A1(new_n75), .A2(new_n644), .ZN(new_n746));
  NOR2_X1   g0682(.A1(new_n76), .A2(new_n552), .ZN(new_n747));
  NOR2_X1   g0683(.A1(new_n89), .A2(new_n468), .ZN(new_n748));
  NOR2_X1   g0684(.A1(new_n110), .A2(new_n392), .ZN(new_n749));
  NOR2_X1   g0685(.A1(new_n139), .A2(new_n324), .ZN(new_n750));
  NOR2_X1   g0686(.A1(new_n176), .A2(new_n264), .ZN(new_n751));
  NOR2_X1   g0687(.A1(new_n221), .A2(new_n212), .ZN(new_n752));
  NOR2_X1   g0688(.A1(new_n274), .A2(new_n168), .ZN(new_n753));
  NOR2_X1   g0689(.A1(new_n335), .A2(new_n132), .ZN(new_n754));
  NOR2_X1   g0690(.A1(new_n404), .A2(new_n104), .ZN(new_n755));
  NOR2_X1   g0691(.A1(new_n481), .A2(new_n84), .ZN(new_n756));
  NOR2_X1   g0692(.A1(new_n566), .A2(new_n72), .ZN(new_n757));
  INV_X1    g0693(.A(new_n660), .ZN(new_n758));
  AOI22_X1  g0694(.A1(G14), .A2(G18), .B1(G15), .B2(G17), .ZN(new_n759));
  INV_X1    g0695(.A(G15), .ZN(new_n760));
  NOR2_X1   g0696(.A1(new_n760), .A2(new_n77), .ZN(new_n761));
  INV_X1    g0697(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g0698(.A1(new_n659), .A2(new_n66), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g0699(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0700(.A(new_n764), .B1(new_n758), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g0701(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0702(.A(new_n766), .B1(new_n757), .B2(new_n765), .ZN(new_n767));
  INV_X1    g0703(.A(new_n767), .ZN(new_n768));
  INV_X1    g0704(.A(new_n661), .ZN(new_n769));
  NOR2_X1   g0705(.A1(new_n769), .A2(new_n663), .ZN(new_n770));
  NOR2_X1   g0706(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0707(.A(new_n771), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  INV_X1    g0708(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0709(.A1(new_n756), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0710(.A(new_n774), .B1(new_n756), .B2(new_n773), .ZN(new_n775));
  INV_X1    g0711(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0712(.A1(new_n668), .A2(new_n671), .ZN(new_n777));
  NOR2_X1   g0713(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0714(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  INV_X1    g0715(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0716(.A1(new_n755), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0717(.A(new_n781), .B1(new_n755), .B2(new_n780), .ZN(new_n782));
  INV_X1    g0718(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0719(.A1(new_n675), .A2(new_n678), .ZN(new_n784));
  NOR2_X1   g0720(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0721(.A(new_n785), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  INV_X1    g0722(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0723(.A1(new_n754), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0724(.A(new_n788), .B1(new_n754), .B2(new_n787), .ZN(new_n789));
  INV_X1    g0725(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0726(.A1(new_n682), .A2(new_n685), .ZN(new_n791));
  NOR2_X1   g0727(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0728(.A(new_n792), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  INV_X1    g0729(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0730(.A1(new_n753), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0731(.A(new_n795), .B1(new_n753), .B2(new_n794), .ZN(new_n796));
  INV_X1    g0732(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0733(.A1(new_n689), .A2(new_n692), .ZN(new_n798));
  NOR2_X1   g0734(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0735(.A(new_n799), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  INV_X1    g0736(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0737(.A1(new_n752), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0738(.A(new_n802), .B1(new_n752), .B2(new_n801), .ZN(new_n803));
  INV_X1    g0739(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0740(.A1(new_n696), .A2(new_n699), .ZN(new_n805));
  NOR2_X1   g0741(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0742(.A(new_n806), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  INV_X1    g0743(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0744(.A1(new_n751), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0745(.A(new_n809), .B1(new_n751), .B2(new_n808), .ZN(new_n810));
  INV_X1    g0746(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0747(.A1(new_n703), .A2(new_n706), .ZN(new_n812));
  NOR2_X1   g0748(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0749(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0750(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0751(.A1(new_n750), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0752(.A(new_n816), .B1(new_n750), .B2(new_n815), .ZN(new_n817));
  INV_X1    g0753(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0754(.A1(new_n710), .A2(new_n713), .ZN(new_n819));
  NOR2_X1   g0755(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0756(.A(new_n820), .B1(new_n818), .B2(new_n819), .ZN(new_n821));
  INV_X1    g0757(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0758(.A1(new_n749), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0759(.A(new_n823), .B1(new_n749), .B2(new_n822), .ZN(new_n824));
  INV_X1    g0760(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0761(.A1(new_n717), .A2(new_n720), .ZN(new_n826));
  NOR2_X1   g0762(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0763(.A(new_n827), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  INV_X1    g0764(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0765(.A1(new_n748), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0766(.A(new_n830), .B1(new_n748), .B2(new_n829), .ZN(new_n831));
  INV_X1    g0767(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0768(.A1(new_n724), .A2(new_n727), .ZN(new_n833));
  NOR2_X1   g0769(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0770(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  INV_X1    g0771(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0772(.A1(new_n747), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0773(.A(new_n837), .B1(new_n747), .B2(new_n836), .ZN(new_n838));
  INV_X1    g0774(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0775(.A1(new_n731), .A2(new_n734), .ZN(new_n840));
  NOR2_X1   g0776(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0777(.A(new_n841), .B1(new_n839), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0778(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0779(.A1(new_n746), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0780(.A(new_n844), .B1(new_n746), .B2(new_n843), .ZN(new_n845));
  INV_X1    g0781(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0782(.A1(new_n738), .A2(new_n741), .ZN(new_n847));
  NOR2_X1   g0783(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0784(.A(new_n848), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  INV_X1    g0785(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0786(.A1(new_n745), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0787(.A(new_n851), .B1(new_n745), .B2(new_n850), .ZN(new_n852));
  INV_X1    g0788(.A(new_n852), .ZN(G6271));
  INV_X1    g0789(.A(G32), .ZN(new_n854));
  NOR2_X1   g0790(.A1(new_n65), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0791(.A1(new_n75), .A2(new_n744), .ZN(new_n856));
  NOR2_X1   g0792(.A1(new_n76), .A2(new_n644), .ZN(new_n857));
  NOR2_X1   g0793(.A1(new_n89), .A2(new_n552), .ZN(new_n858));
  NOR2_X1   g0794(.A1(new_n110), .A2(new_n468), .ZN(new_n859));
  NOR2_X1   g0795(.A1(new_n139), .A2(new_n392), .ZN(new_n860));
  NOR2_X1   g0796(.A1(new_n176), .A2(new_n324), .ZN(new_n861));
  NOR2_X1   g0797(.A1(new_n221), .A2(new_n264), .ZN(new_n862));
  NOR2_X1   g0798(.A1(new_n274), .A2(new_n212), .ZN(new_n863));
  NOR2_X1   g0799(.A1(new_n335), .A2(new_n168), .ZN(new_n864));
  NOR2_X1   g0800(.A1(new_n404), .A2(new_n132), .ZN(new_n865));
  NOR2_X1   g0801(.A1(new_n481), .A2(new_n104), .ZN(new_n866));
  NOR2_X1   g0802(.A1(new_n566), .A2(new_n84), .ZN(new_n867));
  NOR2_X1   g0803(.A1(new_n659), .A2(new_n72), .ZN(new_n868));
  INV_X1    g0804(.A(G16), .ZN(new_n869));
  NOR2_X1   g0805(.A1(new_n869), .A2(new_n66), .ZN(new_n870));
  NAND3_X1  g0806(.A1(new_n659), .A2(new_n761), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g0807(.A(new_n871), .B1(new_n761), .B2(new_n870), .ZN(new_n872));
  AOI21_X1  g0808(.A(new_n872), .B1(new_n869), .B2(new_n763), .ZN(new_n873));
  INV_X1    g0809(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g0810(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0811(.A(new_n875), .B1(new_n868), .B2(new_n874), .ZN(new_n876));
  INV_X1    g0812(.A(new_n876), .ZN(new_n877));
  INV_X1    g0813(.A(new_n764), .ZN(new_n878));
  NOR2_X1   g0814(.A1(new_n878), .A2(new_n766), .ZN(new_n879));
  NOR2_X1   g0815(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0816(.A(new_n880), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  INV_X1    g0817(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g0818(.A1(new_n867), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0819(.A(new_n883), .B1(new_n867), .B2(new_n882), .ZN(new_n884));
  INV_X1    g0820(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g0821(.A1(new_n771), .A2(new_n774), .ZN(new_n886));
  NOR2_X1   g0822(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0823(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  INV_X1    g0824(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g0825(.A1(new_n866), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0826(.A(new_n890), .B1(new_n866), .B2(new_n889), .ZN(new_n891));
  INV_X1    g0827(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0828(.A1(new_n778), .A2(new_n781), .ZN(new_n893));
  NOR2_X1   g0829(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0830(.A(new_n894), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  INV_X1    g0831(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g0832(.A1(new_n865), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0833(.A(new_n897), .B1(new_n865), .B2(new_n896), .ZN(new_n898));
  INV_X1    g0834(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0835(.A1(new_n785), .A2(new_n788), .ZN(new_n900));
  NOR2_X1   g0836(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0837(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  INV_X1    g0838(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g0839(.A1(new_n864), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0840(.A(new_n904), .B1(new_n864), .B2(new_n903), .ZN(new_n905));
  INV_X1    g0841(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0842(.A1(new_n792), .A2(new_n795), .ZN(new_n907));
  NOR2_X1   g0843(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0844(.A(new_n908), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  INV_X1    g0845(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0846(.A1(new_n863), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0847(.A(new_n911), .B1(new_n863), .B2(new_n910), .ZN(new_n912));
  INV_X1    g0848(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0849(.A1(new_n799), .A2(new_n802), .ZN(new_n914));
  NOR2_X1   g0850(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0851(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  INV_X1    g0852(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g0853(.A1(new_n862), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0854(.A(new_n918), .B1(new_n862), .B2(new_n917), .ZN(new_n919));
  INV_X1    g0855(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0856(.A1(new_n806), .A2(new_n809), .ZN(new_n921));
  NOR2_X1   g0857(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0858(.A(new_n922), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  INV_X1    g0859(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0860(.A1(new_n861), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0861(.A(new_n925), .B1(new_n861), .B2(new_n924), .ZN(new_n926));
  INV_X1    g0862(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0863(.A1(new_n813), .A2(new_n816), .ZN(new_n928));
  NOR2_X1   g0864(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0865(.A(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  INV_X1    g0866(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0867(.A1(new_n860), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0868(.A(new_n932), .B1(new_n860), .B2(new_n931), .ZN(new_n933));
  INV_X1    g0869(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0870(.A1(new_n820), .A2(new_n823), .ZN(new_n935));
  NOR2_X1   g0871(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0872(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  INV_X1    g0873(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0874(.A1(new_n859), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0875(.A(new_n939), .B1(new_n859), .B2(new_n938), .ZN(new_n940));
  INV_X1    g0876(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g0877(.A1(new_n827), .A2(new_n830), .ZN(new_n942));
  NOR2_X1   g0878(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0879(.A(new_n943), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  INV_X1    g0880(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0881(.A1(new_n858), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0882(.A(new_n946), .B1(new_n858), .B2(new_n945), .ZN(new_n947));
  INV_X1    g0883(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g0884(.A1(new_n834), .A2(new_n837), .ZN(new_n949));
  NOR2_X1   g0885(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0886(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  INV_X1    g0887(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0888(.A1(new_n857), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0889(.A(new_n953), .B1(new_n857), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0890(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0891(.A1(new_n841), .A2(new_n844), .ZN(new_n956));
  NOR2_X1   g0892(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0893(.A(new_n957), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  INV_X1    g0894(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0895(.A1(new_n856), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0896(.A(new_n960), .B1(new_n856), .B2(new_n959), .ZN(new_n961));
  INV_X1    g0897(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0898(.A1(new_n848), .A2(new_n851), .ZN(new_n963));
  NOR2_X1   g0899(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0900(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0901(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0902(.A1(new_n855), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0903(.A(new_n967), .B1(new_n855), .B2(new_n966), .ZN(new_n968));
  INV_X1    g0904(.A(new_n968), .ZN(G6272));
  NOR2_X1   g0905(.A1(new_n964), .A2(new_n967), .ZN(new_n970));
  NOR2_X1   g0906(.A1(new_n75), .A2(new_n854), .ZN(new_n971));
  NOR2_X1   g0907(.A1(new_n957), .A2(new_n960), .ZN(new_n972));
  NOR2_X1   g0908(.A1(new_n76), .A2(new_n744), .ZN(new_n973));
  NOR2_X1   g0909(.A1(new_n950), .A2(new_n953), .ZN(new_n974));
  NOR2_X1   g0910(.A1(new_n89), .A2(new_n644), .ZN(new_n975));
  NOR2_X1   g0911(.A1(new_n943), .A2(new_n946), .ZN(new_n976));
  NOR2_X1   g0912(.A1(new_n110), .A2(new_n552), .ZN(new_n977));
  NOR2_X1   g0913(.A1(new_n936), .A2(new_n939), .ZN(new_n978));
  NOR2_X1   g0914(.A1(new_n139), .A2(new_n468), .ZN(new_n979));
  NOR2_X1   g0915(.A1(new_n929), .A2(new_n932), .ZN(new_n980));
  NOR2_X1   g0916(.A1(new_n176), .A2(new_n392), .ZN(new_n981));
  NOR2_X1   g0917(.A1(new_n922), .A2(new_n925), .ZN(new_n982));
  NOR2_X1   g0918(.A1(new_n221), .A2(new_n324), .ZN(new_n983));
  NOR2_X1   g0919(.A1(new_n915), .A2(new_n918), .ZN(new_n984));
  NOR2_X1   g0920(.A1(new_n274), .A2(new_n264), .ZN(new_n985));
  NOR2_X1   g0921(.A1(new_n908), .A2(new_n911), .ZN(new_n986));
  NOR2_X1   g0922(.A1(new_n335), .A2(new_n212), .ZN(new_n987));
  NOR2_X1   g0923(.A1(new_n901), .A2(new_n904), .ZN(new_n988));
  NOR2_X1   g0924(.A1(new_n404), .A2(new_n168), .ZN(new_n989));
  NOR2_X1   g0925(.A1(new_n894), .A2(new_n897), .ZN(new_n990));
  NOR2_X1   g0926(.A1(new_n481), .A2(new_n132), .ZN(new_n991));
  NOR2_X1   g0927(.A1(new_n887), .A2(new_n890), .ZN(new_n992));
  NOR2_X1   g0928(.A1(new_n566), .A2(new_n104), .ZN(new_n993));
  NOR2_X1   g0929(.A1(new_n880), .A2(new_n883), .ZN(new_n994));
  NOR2_X1   g0930(.A1(new_n659), .A2(new_n84), .ZN(new_n995));
  NOR2_X1   g0931(.A1(new_n872), .A2(new_n875), .ZN(new_n996));
  NOR2_X1   g0932(.A1(new_n760), .A2(new_n72), .ZN(new_n997));
  OAI211_X1 g0933(.A(G16), .B(G18), .C1(new_n760), .C2(new_n66), .ZN(new_n998));
  XNOR2_X1  g0934(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NOR2_X1   g0935(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0936(.A(new_n1000), .B1(new_n996), .B2(new_n999), .ZN(new_n1001));
  INV_X1    g0937(.A(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0938(.A1(new_n995), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0939(.A(new_n1003), .B1(new_n995), .B2(new_n1002), .ZN(new_n1004));
  INV_X1    g0940(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0941(.A1(new_n994), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0942(.A(new_n1006), .B1(new_n994), .B2(new_n1005), .ZN(new_n1007));
  INV_X1    g0943(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0944(.A1(new_n993), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0945(.A(new_n1009), .B1(new_n993), .B2(new_n1008), .ZN(new_n1010));
  INV_X1    g0946(.A(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0947(.A1(new_n992), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0948(.A(new_n1012), .B1(new_n992), .B2(new_n1011), .ZN(new_n1013));
  INV_X1    g0949(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0950(.A1(new_n991), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0951(.A(new_n1015), .B1(new_n991), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g0952(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0953(.A1(new_n990), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0954(.A(new_n1018), .B1(new_n990), .B2(new_n1017), .ZN(new_n1019));
  INV_X1    g0955(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0956(.A1(new_n989), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0957(.A(new_n1021), .B1(new_n989), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g0958(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0959(.A1(new_n988), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0960(.A(new_n1024), .B1(new_n988), .B2(new_n1023), .ZN(new_n1025));
  INV_X1    g0961(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0962(.A1(new_n987), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0963(.A(new_n1027), .B1(new_n987), .B2(new_n1026), .ZN(new_n1028));
  INV_X1    g0964(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0965(.A1(new_n986), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0966(.A(new_n1030), .B1(new_n986), .B2(new_n1029), .ZN(new_n1031));
  INV_X1    g0967(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0968(.A1(new_n985), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0969(.A(new_n1033), .B1(new_n985), .B2(new_n1032), .ZN(new_n1034));
  INV_X1    g0970(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0971(.A1(new_n984), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0972(.A(new_n1036), .B1(new_n984), .B2(new_n1035), .ZN(new_n1037));
  INV_X1    g0973(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0974(.A1(new_n983), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0975(.A(new_n1039), .B1(new_n983), .B2(new_n1038), .ZN(new_n1040));
  INV_X1    g0976(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0977(.A1(new_n982), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0978(.A(new_n1042), .B1(new_n982), .B2(new_n1041), .ZN(new_n1043));
  INV_X1    g0979(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0980(.A1(new_n981), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0981(.A(new_n1045), .B1(new_n981), .B2(new_n1044), .ZN(new_n1046));
  INV_X1    g0982(.A(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0983(.A1(new_n980), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0984(.A(new_n1048), .B1(new_n980), .B2(new_n1047), .ZN(new_n1049));
  INV_X1    g0985(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0986(.A1(new_n979), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0987(.A(new_n1051), .B1(new_n979), .B2(new_n1050), .ZN(new_n1052));
  INV_X1    g0988(.A(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0989(.A1(new_n978), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0990(.A(new_n1054), .B1(new_n978), .B2(new_n1053), .ZN(new_n1055));
  INV_X1    g0991(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0992(.A1(new_n977), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0993(.A(new_n1057), .B1(new_n977), .B2(new_n1056), .ZN(new_n1058));
  INV_X1    g0994(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0995(.A1(new_n976), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0996(.A(new_n1060), .B1(new_n976), .B2(new_n1059), .ZN(new_n1061));
  INV_X1    g0997(.A(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0998(.A1(new_n975), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0999(.A(new_n1063), .B1(new_n975), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g1000(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g1001(.A1(new_n974), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g1002(.A(new_n1066), .B1(new_n974), .B2(new_n1065), .ZN(new_n1067));
  INV_X1    g1003(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g1004(.A1(new_n973), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g1005(.A(new_n1069), .B1(new_n973), .B2(new_n1068), .ZN(new_n1070));
  INV_X1    g1006(.A(new_n1070), .ZN(new_n1071));
  NOR2_X1   g1007(.A1(new_n972), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g1008(.A(new_n1072), .B1(new_n972), .B2(new_n1071), .ZN(new_n1073));
  INV_X1    g1009(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g1010(.A1(new_n971), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g1011(.A(new_n1075), .B1(new_n971), .B2(new_n1074), .ZN(new_n1076));
  INV_X1    g1012(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g1013(.A1(new_n970), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g1014(.A(new_n1078), .B1(new_n970), .B2(new_n1077), .ZN(new_n1079));
  INV_X1    g1015(.A(new_n1079), .ZN(G6273));
  NOR2_X1   g1016(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1081));
  NOR2_X1   g1017(.A1(new_n76), .A2(new_n854), .ZN(new_n1082));
  NOR2_X1   g1018(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1083));
  NOR2_X1   g1019(.A1(new_n89), .A2(new_n744), .ZN(new_n1084));
  NOR2_X1   g1020(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1085));
  NOR2_X1   g1021(.A1(new_n110), .A2(new_n644), .ZN(new_n1086));
  NOR2_X1   g1022(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1087));
  NOR2_X1   g1023(.A1(new_n139), .A2(new_n552), .ZN(new_n1088));
  NOR2_X1   g1024(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1089));
  NOR2_X1   g1025(.A1(new_n176), .A2(new_n468), .ZN(new_n1090));
  NOR2_X1   g1026(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1091));
  NOR2_X1   g1027(.A1(new_n221), .A2(new_n392), .ZN(new_n1092));
  NOR2_X1   g1028(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1093));
  NOR2_X1   g1029(.A1(new_n274), .A2(new_n324), .ZN(new_n1094));
  NOR2_X1   g1030(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1095));
  NOR2_X1   g1031(.A1(new_n335), .A2(new_n264), .ZN(new_n1096));
  NOR2_X1   g1032(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1097));
  NOR2_X1   g1033(.A1(new_n404), .A2(new_n212), .ZN(new_n1098));
  NOR2_X1   g1034(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1099));
  NOR2_X1   g1035(.A1(new_n481), .A2(new_n168), .ZN(new_n1100));
  NOR2_X1   g1036(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1101));
  NOR2_X1   g1037(.A1(new_n566), .A2(new_n132), .ZN(new_n1102));
  NOR2_X1   g1038(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1103));
  NOR2_X1   g1039(.A1(new_n659), .A2(new_n104), .ZN(new_n1104));
  NOR2_X1   g1040(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1105));
  NOR2_X1   g1041(.A1(new_n760), .A2(new_n84), .ZN(new_n1106));
  NOR2_X1   g1042(.A1(new_n66), .A2(new_n762), .ZN(new_n1107));
  OAI21_X1  g1043(.A(G16), .B1(G19), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g1044(.A(new_n1108), .B1(G18), .B2(new_n997), .ZN(new_n1109));
  INV_X1    g1045(.A(new_n1109), .ZN(new_n1110));
  NOR2_X1   g1046(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g1047(.A(new_n1111), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1112));
  INV_X1    g1048(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g1049(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g1050(.A(new_n1114), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1115));
  INV_X1    g1051(.A(new_n1115), .ZN(new_n1116));
  NOR2_X1   g1052(.A1(new_n1104), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g1053(.A(new_n1117), .B1(new_n1104), .B2(new_n1116), .ZN(new_n1118));
  INV_X1    g1054(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g1055(.A1(new_n1103), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g1056(.A(new_n1120), .B1(new_n1103), .B2(new_n1119), .ZN(new_n1121));
  INV_X1    g1057(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g1058(.A1(new_n1102), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g1059(.A(new_n1123), .B1(new_n1102), .B2(new_n1122), .ZN(new_n1124));
  INV_X1    g1060(.A(new_n1124), .ZN(new_n1125));
  NOR2_X1   g1061(.A1(new_n1101), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g1062(.A(new_n1126), .B1(new_n1101), .B2(new_n1125), .ZN(new_n1127));
  INV_X1    g1063(.A(new_n1127), .ZN(new_n1128));
  NOR2_X1   g1064(.A1(new_n1100), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g1065(.A(new_n1129), .B1(new_n1100), .B2(new_n1128), .ZN(new_n1130));
  INV_X1    g1066(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g1067(.A1(new_n1099), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g1068(.A(new_n1132), .B1(new_n1099), .B2(new_n1131), .ZN(new_n1133));
  INV_X1    g1069(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g1070(.A1(new_n1098), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g1071(.A(new_n1135), .B1(new_n1098), .B2(new_n1134), .ZN(new_n1136));
  INV_X1    g1072(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g1073(.A1(new_n1097), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g1074(.A(new_n1138), .B1(new_n1097), .B2(new_n1137), .ZN(new_n1139));
  INV_X1    g1075(.A(new_n1139), .ZN(new_n1140));
  NOR2_X1   g1076(.A1(new_n1096), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g1077(.A(new_n1141), .B1(new_n1096), .B2(new_n1140), .ZN(new_n1142));
  INV_X1    g1078(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g1079(.A1(new_n1095), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g1080(.A(new_n1144), .B1(new_n1095), .B2(new_n1143), .ZN(new_n1145));
  INV_X1    g1081(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g1082(.A1(new_n1094), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g1083(.A(new_n1147), .B1(new_n1094), .B2(new_n1146), .ZN(new_n1148));
  INV_X1    g1084(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g1085(.A1(new_n1093), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g1086(.A(new_n1150), .B1(new_n1093), .B2(new_n1149), .ZN(new_n1151));
  INV_X1    g1087(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g1088(.A1(new_n1092), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g1089(.A(new_n1153), .B1(new_n1092), .B2(new_n1152), .ZN(new_n1154));
  INV_X1    g1090(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g1091(.A1(new_n1091), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g1092(.A(new_n1156), .B1(new_n1091), .B2(new_n1155), .ZN(new_n1157));
  INV_X1    g1093(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g1094(.A1(new_n1090), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g1095(.A(new_n1159), .B1(new_n1090), .B2(new_n1158), .ZN(new_n1160));
  INV_X1    g1096(.A(new_n1160), .ZN(new_n1161));
  NOR2_X1   g1097(.A1(new_n1089), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g1098(.A(new_n1162), .B1(new_n1089), .B2(new_n1161), .ZN(new_n1163));
  INV_X1    g1099(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g1100(.A1(new_n1088), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g1101(.A(new_n1165), .B1(new_n1088), .B2(new_n1164), .ZN(new_n1166));
  INV_X1    g1102(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g1103(.A1(new_n1087), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g1104(.A(new_n1168), .B1(new_n1087), .B2(new_n1167), .ZN(new_n1169));
  INV_X1    g1105(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g1106(.A1(new_n1086), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g1107(.A(new_n1171), .B1(new_n1086), .B2(new_n1170), .ZN(new_n1172));
  INV_X1    g1108(.A(new_n1172), .ZN(new_n1173));
  NOR2_X1   g1109(.A1(new_n1085), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g1110(.A(new_n1174), .B1(new_n1085), .B2(new_n1173), .ZN(new_n1175));
  INV_X1    g1111(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g1112(.A1(new_n1084), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g1113(.A(new_n1177), .B1(new_n1084), .B2(new_n1176), .ZN(new_n1178));
  INV_X1    g1114(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g1115(.A1(new_n1083), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g1116(.A(new_n1180), .B1(new_n1083), .B2(new_n1179), .ZN(new_n1181));
  INV_X1    g1117(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g1118(.A1(new_n1082), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g1119(.A(new_n1183), .B1(new_n1082), .B2(new_n1182), .ZN(new_n1184));
  INV_X1    g1120(.A(new_n1184), .ZN(new_n1185));
  NOR2_X1   g1121(.A1(new_n1081), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g1122(.A(new_n1186), .B1(new_n1081), .B2(new_n1185), .ZN(new_n1187));
  XNOR2_X1  g1123(.A(new_n1078), .B(new_n1187), .ZN(G6274));
  AOI21_X1  g1124(.A(new_n1186), .B1(new_n1078), .B2(new_n1187), .ZN(new_n1189));
  NOR2_X1   g1125(.A1(new_n89), .A2(new_n854), .ZN(new_n1190));
  NOR2_X1   g1126(.A1(new_n110), .A2(new_n744), .ZN(new_n1191));
  NOR2_X1   g1127(.A1(new_n139), .A2(new_n644), .ZN(new_n1192));
  NOR2_X1   g1128(.A1(new_n176), .A2(new_n552), .ZN(new_n1193));
  NOR2_X1   g1129(.A1(new_n221), .A2(new_n468), .ZN(new_n1194));
  NOR2_X1   g1130(.A1(new_n274), .A2(new_n392), .ZN(new_n1195));
  NOR2_X1   g1131(.A1(new_n335), .A2(new_n324), .ZN(new_n1196));
  NOR2_X1   g1132(.A1(new_n404), .A2(new_n264), .ZN(new_n1197));
  NOR2_X1   g1133(.A1(new_n481), .A2(new_n212), .ZN(new_n1198));
  NOR2_X1   g1134(.A1(new_n566), .A2(new_n168), .ZN(new_n1199));
  NOR2_X1   g1135(.A1(new_n659), .A2(new_n132), .ZN(new_n1200));
  NOR2_X1   g1136(.A1(new_n760), .A2(new_n104), .ZN(new_n1201));
  OR2_X1    g1137(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1202));
  OAI21_X1  g1138(.A(new_n1202), .B1(new_n869), .B2(new_n84), .ZN(new_n1203));
  OAI21_X1  g1139(.A(new_n1203), .B1(new_n84), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1140(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1141(.A(new_n1205), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1206));
  INV_X1    g1142(.A(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1143(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1208));
  NOR2_X1   g1144(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1145(.A(new_n1209), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1210));
  INV_X1    g1146(.A(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1147(.A1(new_n1200), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1148(.A(new_n1212), .B1(new_n1200), .B2(new_n1211), .ZN(new_n1213));
  INV_X1    g1149(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1150(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1215));
  NOR2_X1   g1151(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1152(.A(new_n1216), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1217));
  INV_X1    g1153(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1154(.A1(new_n1199), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1155(.A(new_n1219), .B1(new_n1199), .B2(new_n1218), .ZN(new_n1220));
  INV_X1    g1156(.A(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1157(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1222));
  NOR2_X1   g1158(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1159(.A(new_n1223), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1224));
  INV_X1    g1160(.A(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1161(.A1(new_n1198), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1162(.A(new_n1226), .B1(new_n1198), .B2(new_n1225), .ZN(new_n1227));
  INV_X1    g1163(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1164(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1229));
  NOR2_X1   g1165(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1166(.A(new_n1230), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1231));
  INV_X1    g1167(.A(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1168(.A1(new_n1197), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1169(.A(new_n1233), .B1(new_n1197), .B2(new_n1232), .ZN(new_n1234));
  INV_X1    g1170(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1171(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1236));
  NOR2_X1   g1172(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1173(.A(new_n1237), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1238));
  INV_X1    g1174(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1175(.A1(new_n1196), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1176(.A(new_n1240), .B1(new_n1196), .B2(new_n1239), .ZN(new_n1241));
  INV_X1    g1177(.A(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1178(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1243));
  NOR2_X1   g1179(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1180(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1245));
  INV_X1    g1181(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1182(.A1(new_n1195), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1183(.A(new_n1247), .B1(new_n1195), .B2(new_n1246), .ZN(new_n1248));
  INV_X1    g1184(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1185(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1250));
  NOR2_X1   g1186(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1187(.A(new_n1251), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1252));
  INV_X1    g1188(.A(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1189(.A1(new_n1194), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1190(.A(new_n1254), .B1(new_n1194), .B2(new_n1253), .ZN(new_n1255));
  INV_X1    g1191(.A(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1192(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1257));
  NOR2_X1   g1193(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1194(.A(new_n1258), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1259));
  INV_X1    g1195(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1196(.A1(new_n1193), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1197(.A(new_n1261), .B1(new_n1193), .B2(new_n1260), .ZN(new_n1262));
  INV_X1    g1198(.A(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1199(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1264));
  NOR2_X1   g1200(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1201(.A(new_n1265), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1266));
  INV_X1    g1202(.A(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1203(.A1(new_n1192), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1204(.A(new_n1268), .B1(new_n1192), .B2(new_n1267), .ZN(new_n1269));
  INV_X1    g1205(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1206(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1271));
  NOR2_X1   g1207(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1208(.A(new_n1272), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1273));
  INV_X1    g1209(.A(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1210(.A1(new_n1191), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1211(.A(new_n1275), .B1(new_n1191), .B2(new_n1274), .ZN(new_n1276));
  INV_X1    g1212(.A(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1213(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1278));
  NOR2_X1   g1214(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1215(.A(new_n1279), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1280));
  INV_X1    g1216(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1217(.A1(new_n1190), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1218(.A(new_n1282), .B1(new_n1190), .B2(new_n1281), .ZN(new_n1283));
  INV_X1    g1219(.A(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1220(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1285));
  NOR2_X1   g1221(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1222(.A(new_n1286), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1287));
  INV_X1    g1223(.A(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1224(.A1(new_n1189), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1225(.A(new_n1289), .B1(new_n1189), .B2(new_n1288), .ZN(new_n1290));
  INV_X1    g1226(.A(new_n1290), .ZN(G6275));
  NOR2_X1   g1227(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1292));
  NOR2_X1   g1228(.A1(new_n110), .A2(new_n854), .ZN(new_n1293));
  NOR2_X1   g1229(.A1(new_n139), .A2(new_n744), .ZN(new_n1294));
  NOR2_X1   g1230(.A1(new_n176), .A2(new_n644), .ZN(new_n1295));
  NOR2_X1   g1231(.A1(new_n221), .A2(new_n552), .ZN(new_n1296));
  NOR2_X1   g1232(.A1(new_n274), .A2(new_n468), .ZN(new_n1297));
  NOR2_X1   g1233(.A1(new_n335), .A2(new_n392), .ZN(new_n1298));
  NOR2_X1   g1234(.A1(new_n404), .A2(new_n324), .ZN(new_n1299));
  NOR2_X1   g1235(.A1(new_n481), .A2(new_n264), .ZN(new_n1300));
  NOR2_X1   g1236(.A1(new_n566), .A2(new_n212), .ZN(new_n1301));
  NOR2_X1   g1237(.A1(new_n659), .A2(new_n168), .ZN(new_n1302));
  NOR2_X1   g1238(.A1(new_n760), .A2(new_n132), .ZN(new_n1303));
  NOR2_X1   g1239(.A1(new_n869), .A2(new_n104), .ZN(new_n1304));
  INV_X1    g1240(.A(new_n1203), .ZN(new_n1305));
  NOR2_X1   g1241(.A1(new_n1305), .A2(new_n1205), .ZN(new_n1306));
  NOR2_X1   g1242(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1243(.A(new_n1307), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1308));
  INV_X1    g1244(.A(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1245(.A1(new_n1303), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1246(.A(new_n1310), .B1(new_n1303), .B2(new_n1309), .ZN(new_n1311));
  INV_X1    g1247(.A(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1248(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1313));
  NOR2_X1   g1249(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1250(.A(new_n1314), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1315));
  INV_X1    g1251(.A(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1252(.A1(new_n1302), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1253(.A(new_n1317), .B1(new_n1302), .B2(new_n1316), .ZN(new_n1318));
  INV_X1    g1254(.A(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1255(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1320));
  NOR2_X1   g1256(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1257(.A(new_n1321), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1322));
  INV_X1    g1258(.A(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1259(.A1(new_n1301), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1260(.A(new_n1324), .B1(new_n1301), .B2(new_n1323), .ZN(new_n1325));
  INV_X1    g1261(.A(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1262(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1327));
  NOR2_X1   g1263(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1264(.A(new_n1328), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1329));
  INV_X1    g1265(.A(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1266(.A1(new_n1300), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1267(.A(new_n1331), .B1(new_n1300), .B2(new_n1330), .ZN(new_n1332));
  INV_X1    g1268(.A(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1269(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1334));
  NOR2_X1   g1270(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1271(.A(new_n1335), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1336));
  INV_X1    g1272(.A(new_n1336), .ZN(new_n1337));
  NOR2_X1   g1273(.A1(new_n1299), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1274(.A(new_n1338), .B1(new_n1299), .B2(new_n1337), .ZN(new_n1339));
  INV_X1    g1275(.A(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1276(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1341));
  NOR2_X1   g1277(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1278(.A(new_n1342), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1343));
  INV_X1    g1279(.A(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1280(.A1(new_n1298), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1281(.A(new_n1345), .B1(new_n1298), .B2(new_n1344), .ZN(new_n1346));
  INV_X1    g1282(.A(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1283(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1348));
  NOR2_X1   g1284(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1285(.A(new_n1349), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1350));
  INV_X1    g1286(.A(new_n1350), .ZN(new_n1351));
  NOR2_X1   g1287(.A1(new_n1297), .A2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1288(.A(new_n1352), .B1(new_n1297), .B2(new_n1351), .ZN(new_n1353));
  INV_X1    g1289(.A(new_n1353), .ZN(new_n1354));
  NOR2_X1   g1290(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1355));
  NOR2_X1   g1291(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1292(.A(new_n1356), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1357));
  INV_X1    g1293(.A(new_n1357), .ZN(new_n1358));
  NOR2_X1   g1294(.A1(new_n1296), .A2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1295(.A(new_n1359), .B1(new_n1296), .B2(new_n1358), .ZN(new_n1360));
  INV_X1    g1296(.A(new_n1360), .ZN(new_n1361));
  NOR2_X1   g1297(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1362));
  NOR2_X1   g1298(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1299(.A(new_n1363), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1364));
  INV_X1    g1300(.A(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1301(.A1(new_n1295), .A2(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1302(.A(new_n1366), .B1(new_n1295), .B2(new_n1365), .ZN(new_n1367));
  INV_X1    g1303(.A(new_n1367), .ZN(new_n1368));
  NOR2_X1   g1304(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1369));
  NOR2_X1   g1305(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1306(.A(new_n1370), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1371));
  INV_X1    g1307(.A(new_n1371), .ZN(new_n1372));
  NOR2_X1   g1308(.A1(new_n1294), .A2(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1309(.A(new_n1373), .B1(new_n1294), .B2(new_n1372), .ZN(new_n1374));
  INV_X1    g1310(.A(new_n1374), .ZN(new_n1375));
  NOR2_X1   g1311(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1376));
  NOR2_X1   g1312(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1313(.A(new_n1377), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1378));
  INV_X1    g1314(.A(new_n1378), .ZN(new_n1379));
  NOR2_X1   g1315(.A1(new_n1293), .A2(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1316(.A(new_n1380), .B1(new_n1293), .B2(new_n1379), .ZN(new_n1381));
  INV_X1    g1317(.A(new_n1381), .ZN(new_n1382));
  NOR2_X1   g1318(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1383));
  NOR2_X1   g1319(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1320(.A(new_n1384), .B1(new_n1382), .B2(new_n1383), .ZN(new_n1385));
  INV_X1    g1321(.A(new_n1385), .ZN(new_n1386));
  NOR2_X1   g1322(.A1(new_n1292), .A2(new_n1386), .ZN(new_n1387));
  AOI21_X1  g1323(.A(new_n1387), .B1(new_n1292), .B2(new_n1386), .ZN(new_n1388));
  INV_X1    g1324(.A(new_n1388), .ZN(G6276));
  NOR2_X1   g1325(.A1(new_n1384), .A2(new_n1387), .ZN(new_n1390));
  NOR2_X1   g1326(.A1(new_n139), .A2(new_n854), .ZN(new_n1391));
  NOR2_X1   g1327(.A1(new_n176), .A2(new_n744), .ZN(new_n1392));
  NOR2_X1   g1328(.A1(new_n221), .A2(new_n644), .ZN(new_n1393));
  NOR2_X1   g1329(.A1(new_n274), .A2(new_n552), .ZN(new_n1394));
  NOR2_X1   g1330(.A1(new_n335), .A2(new_n468), .ZN(new_n1395));
  NOR2_X1   g1331(.A1(new_n404), .A2(new_n392), .ZN(new_n1396));
  NOR2_X1   g1332(.A1(new_n481), .A2(new_n324), .ZN(new_n1397));
  NOR2_X1   g1333(.A1(new_n566), .A2(new_n264), .ZN(new_n1398));
  NOR2_X1   g1334(.A1(new_n659), .A2(new_n212), .ZN(new_n1399));
  NOR2_X1   g1335(.A1(new_n760), .A2(new_n168), .ZN(new_n1400));
  NOR2_X1   g1336(.A1(new_n869), .A2(new_n132), .ZN(new_n1401));
  NOR2_X1   g1337(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1402));
  NOR2_X1   g1338(.A1(new_n1401), .A2(new_n1402), .ZN(new_n1403));
  AOI21_X1  g1339(.A(new_n1403), .B1(new_n1401), .B2(new_n1402), .ZN(new_n1404));
  INV_X1    g1340(.A(new_n1404), .ZN(new_n1405));
  NOR2_X1   g1341(.A1(new_n1400), .A2(new_n1405), .ZN(new_n1406));
  AOI21_X1  g1342(.A(new_n1406), .B1(new_n1400), .B2(new_n1405), .ZN(new_n1407));
  INV_X1    g1343(.A(new_n1407), .ZN(new_n1408));
  NOR2_X1   g1344(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1409));
  NOR2_X1   g1345(.A1(new_n1408), .A2(new_n1409), .ZN(new_n1410));
  AOI21_X1  g1346(.A(new_n1410), .B1(new_n1408), .B2(new_n1409), .ZN(new_n1411));
  INV_X1    g1347(.A(new_n1411), .ZN(new_n1412));
  NOR2_X1   g1348(.A1(new_n1399), .A2(new_n1412), .ZN(new_n1413));
  AOI21_X1  g1349(.A(new_n1413), .B1(new_n1399), .B2(new_n1412), .ZN(new_n1414));
  INV_X1    g1350(.A(new_n1414), .ZN(new_n1415));
  NOR2_X1   g1351(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1416));
  NOR2_X1   g1352(.A1(new_n1415), .A2(new_n1416), .ZN(new_n1417));
  AOI21_X1  g1353(.A(new_n1417), .B1(new_n1415), .B2(new_n1416), .ZN(new_n1418));
  INV_X1    g1354(.A(new_n1418), .ZN(new_n1419));
  NOR2_X1   g1355(.A1(new_n1398), .A2(new_n1419), .ZN(new_n1420));
  AOI21_X1  g1356(.A(new_n1420), .B1(new_n1398), .B2(new_n1419), .ZN(new_n1421));
  INV_X1    g1357(.A(new_n1421), .ZN(new_n1422));
  NOR2_X1   g1358(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1423));
  NOR2_X1   g1359(.A1(new_n1422), .A2(new_n1423), .ZN(new_n1424));
  AOI21_X1  g1360(.A(new_n1424), .B1(new_n1422), .B2(new_n1423), .ZN(new_n1425));
  INV_X1    g1361(.A(new_n1425), .ZN(new_n1426));
  NOR2_X1   g1362(.A1(new_n1397), .A2(new_n1426), .ZN(new_n1427));
  AOI21_X1  g1363(.A(new_n1427), .B1(new_n1397), .B2(new_n1426), .ZN(new_n1428));
  INV_X1    g1364(.A(new_n1428), .ZN(new_n1429));
  NOR2_X1   g1365(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1430));
  NOR2_X1   g1366(.A1(new_n1429), .A2(new_n1430), .ZN(new_n1431));
  AOI21_X1  g1367(.A(new_n1431), .B1(new_n1429), .B2(new_n1430), .ZN(new_n1432));
  INV_X1    g1368(.A(new_n1432), .ZN(new_n1433));
  NOR2_X1   g1369(.A1(new_n1396), .A2(new_n1433), .ZN(new_n1434));
  AOI21_X1  g1370(.A(new_n1434), .B1(new_n1396), .B2(new_n1433), .ZN(new_n1435));
  INV_X1    g1371(.A(new_n1435), .ZN(new_n1436));
  NOR2_X1   g1372(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1437));
  NOR2_X1   g1373(.A1(new_n1436), .A2(new_n1437), .ZN(new_n1438));
  AOI21_X1  g1374(.A(new_n1438), .B1(new_n1436), .B2(new_n1437), .ZN(new_n1439));
  INV_X1    g1375(.A(new_n1439), .ZN(new_n1440));
  NOR2_X1   g1376(.A1(new_n1395), .A2(new_n1440), .ZN(new_n1441));
  AOI21_X1  g1377(.A(new_n1441), .B1(new_n1395), .B2(new_n1440), .ZN(new_n1442));
  INV_X1    g1378(.A(new_n1442), .ZN(new_n1443));
  NOR2_X1   g1379(.A1(new_n1349), .A2(new_n1352), .ZN(new_n1444));
  NOR2_X1   g1380(.A1(new_n1443), .A2(new_n1444), .ZN(new_n1445));
  AOI21_X1  g1381(.A(new_n1445), .B1(new_n1443), .B2(new_n1444), .ZN(new_n1446));
  INV_X1    g1382(.A(new_n1446), .ZN(new_n1447));
  NOR2_X1   g1383(.A1(new_n1394), .A2(new_n1447), .ZN(new_n1448));
  AOI21_X1  g1384(.A(new_n1448), .B1(new_n1394), .B2(new_n1447), .ZN(new_n1449));
  INV_X1    g1385(.A(new_n1449), .ZN(new_n1450));
  NOR2_X1   g1386(.A1(new_n1356), .A2(new_n1359), .ZN(new_n1451));
  NOR2_X1   g1387(.A1(new_n1450), .A2(new_n1451), .ZN(new_n1452));
  AOI21_X1  g1388(.A(new_n1452), .B1(new_n1450), .B2(new_n1451), .ZN(new_n1453));
  INV_X1    g1389(.A(new_n1453), .ZN(new_n1454));
  NOR2_X1   g1390(.A1(new_n1393), .A2(new_n1454), .ZN(new_n1455));
  AOI21_X1  g1391(.A(new_n1455), .B1(new_n1393), .B2(new_n1454), .ZN(new_n1456));
  INV_X1    g1392(.A(new_n1456), .ZN(new_n1457));
  NOR2_X1   g1393(.A1(new_n1363), .A2(new_n1366), .ZN(new_n1458));
  NOR2_X1   g1394(.A1(new_n1457), .A2(new_n1458), .ZN(new_n1459));
  AOI21_X1  g1395(.A(new_n1459), .B1(new_n1457), .B2(new_n1458), .ZN(new_n1460));
  INV_X1    g1396(.A(new_n1460), .ZN(new_n1461));
  NOR2_X1   g1397(.A1(new_n1392), .A2(new_n1461), .ZN(new_n1462));
  AOI21_X1  g1398(.A(new_n1462), .B1(new_n1392), .B2(new_n1461), .ZN(new_n1463));
  INV_X1    g1399(.A(new_n1463), .ZN(new_n1464));
  NOR2_X1   g1400(.A1(new_n1370), .A2(new_n1373), .ZN(new_n1465));
  NOR2_X1   g1401(.A1(new_n1464), .A2(new_n1465), .ZN(new_n1466));
  AOI21_X1  g1402(.A(new_n1466), .B1(new_n1464), .B2(new_n1465), .ZN(new_n1467));
  INV_X1    g1403(.A(new_n1467), .ZN(new_n1468));
  NOR2_X1   g1404(.A1(new_n1391), .A2(new_n1468), .ZN(new_n1469));
  AOI21_X1  g1405(.A(new_n1469), .B1(new_n1391), .B2(new_n1468), .ZN(new_n1470));
  INV_X1    g1406(.A(new_n1470), .ZN(new_n1471));
  NOR2_X1   g1407(.A1(new_n1377), .A2(new_n1380), .ZN(new_n1472));
  NOR2_X1   g1408(.A1(new_n1471), .A2(new_n1472), .ZN(new_n1473));
  AOI21_X1  g1409(.A(new_n1473), .B1(new_n1471), .B2(new_n1472), .ZN(new_n1474));
  INV_X1    g1410(.A(new_n1474), .ZN(new_n1475));
  NOR2_X1   g1411(.A1(new_n1390), .A2(new_n1475), .ZN(new_n1476));
  AOI21_X1  g1412(.A(new_n1476), .B1(new_n1390), .B2(new_n1475), .ZN(new_n1477));
  INV_X1    g1413(.A(new_n1477), .ZN(G6277));
  NOR2_X1   g1414(.A1(new_n1473), .A2(new_n1476), .ZN(new_n1479));
  NOR2_X1   g1415(.A1(new_n176), .A2(new_n854), .ZN(new_n1480));
  NOR2_X1   g1416(.A1(new_n221), .A2(new_n744), .ZN(new_n1481));
  NOR2_X1   g1417(.A1(new_n274), .A2(new_n644), .ZN(new_n1482));
  NOR2_X1   g1418(.A1(new_n335), .A2(new_n552), .ZN(new_n1483));
  NOR2_X1   g1419(.A1(new_n404), .A2(new_n468), .ZN(new_n1484));
  NOR2_X1   g1420(.A1(new_n481), .A2(new_n392), .ZN(new_n1485));
  NOR2_X1   g1421(.A1(new_n566), .A2(new_n324), .ZN(new_n1486));
  NOR2_X1   g1422(.A1(new_n659), .A2(new_n264), .ZN(new_n1487));
  NOR2_X1   g1423(.A1(new_n760), .A2(new_n212), .ZN(new_n1488));
  NOR2_X1   g1424(.A1(new_n869), .A2(new_n168), .ZN(new_n1489));
  NOR2_X1   g1425(.A1(new_n1403), .A2(new_n1406), .ZN(new_n1490));
  NOR2_X1   g1426(.A1(new_n1489), .A2(new_n1490), .ZN(new_n1491));
  AOI21_X1  g1427(.A(new_n1491), .B1(new_n1489), .B2(new_n1490), .ZN(new_n1492));
  INV_X1    g1428(.A(new_n1492), .ZN(new_n1493));
  NOR2_X1   g1429(.A1(new_n1488), .A2(new_n1493), .ZN(new_n1494));
  AOI21_X1  g1430(.A(new_n1494), .B1(new_n1488), .B2(new_n1493), .ZN(new_n1495));
  INV_X1    g1431(.A(new_n1495), .ZN(new_n1496));
  NOR2_X1   g1432(.A1(new_n1410), .A2(new_n1413), .ZN(new_n1497));
  NOR2_X1   g1433(.A1(new_n1496), .A2(new_n1497), .ZN(new_n1498));
  AOI21_X1  g1434(.A(new_n1498), .B1(new_n1496), .B2(new_n1497), .ZN(new_n1499));
  INV_X1    g1435(.A(new_n1499), .ZN(new_n1500));
  NOR2_X1   g1436(.A1(new_n1487), .A2(new_n1500), .ZN(new_n1501));
  AOI21_X1  g1437(.A(new_n1501), .B1(new_n1487), .B2(new_n1500), .ZN(new_n1502));
  INV_X1    g1438(.A(new_n1502), .ZN(new_n1503));
  NOR2_X1   g1439(.A1(new_n1417), .A2(new_n1420), .ZN(new_n1504));
  NOR2_X1   g1440(.A1(new_n1503), .A2(new_n1504), .ZN(new_n1505));
  AOI21_X1  g1441(.A(new_n1505), .B1(new_n1503), .B2(new_n1504), .ZN(new_n1506));
  INV_X1    g1442(.A(new_n1506), .ZN(new_n1507));
  NOR2_X1   g1443(.A1(new_n1486), .A2(new_n1507), .ZN(new_n1508));
  AOI21_X1  g1444(.A(new_n1508), .B1(new_n1486), .B2(new_n1507), .ZN(new_n1509));
  INV_X1    g1445(.A(new_n1509), .ZN(new_n1510));
  NOR2_X1   g1446(.A1(new_n1424), .A2(new_n1427), .ZN(new_n1511));
  NOR2_X1   g1447(.A1(new_n1510), .A2(new_n1511), .ZN(new_n1512));
  AOI21_X1  g1448(.A(new_n1512), .B1(new_n1510), .B2(new_n1511), .ZN(new_n1513));
  INV_X1    g1449(.A(new_n1513), .ZN(new_n1514));
  NOR2_X1   g1450(.A1(new_n1485), .A2(new_n1514), .ZN(new_n1515));
  AOI21_X1  g1451(.A(new_n1515), .B1(new_n1485), .B2(new_n1514), .ZN(new_n1516));
  INV_X1    g1452(.A(new_n1516), .ZN(new_n1517));
  NOR2_X1   g1453(.A1(new_n1431), .A2(new_n1434), .ZN(new_n1518));
  NOR2_X1   g1454(.A1(new_n1517), .A2(new_n1518), .ZN(new_n1519));
  AOI21_X1  g1455(.A(new_n1519), .B1(new_n1517), .B2(new_n1518), .ZN(new_n1520));
  INV_X1    g1456(.A(new_n1520), .ZN(new_n1521));
  NOR2_X1   g1457(.A1(new_n1484), .A2(new_n1521), .ZN(new_n1522));
  AOI21_X1  g1458(.A(new_n1522), .B1(new_n1484), .B2(new_n1521), .ZN(new_n1523));
  INV_X1    g1459(.A(new_n1523), .ZN(new_n1524));
  NOR2_X1   g1460(.A1(new_n1438), .A2(new_n1441), .ZN(new_n1525));
  NOR2_X1   g1461(.A1(new_n1524), .A2(new_n1525), .ZN(new_n1526));
  AOI21_X1  g1462(.A(new_n1526), .B1(new_n1524), .B2(new_n1525), .ZN(new_n1527));
  INV_X1    g1463(.A(new_n1527), .ZN(new_n1528));
  NOR2_X1   g1464(.A1(new_n1483), .A2(new_n1528), .ZN(new_n1529));
  AOI21_X1  g1465(.A(new_n1529), .B1(new_n1483), .B2(new_n1528), .ZN(new_n1530));
  INV_X1    g1466(.A(new_n1530), .ZN(new_n1531));
  NOR2_X1   g1467(.A1(new_n1445), .A2(new_n1448), .ZN(new_n1532));
  NOR2_X1   g1468(.A1(new_n1531), .A2(new_n1532), .ZN(new_n1533));
  AOI21_X1  g1469(.A(new_n1533), .B1(new_n1531), .B2(new_n1532), .ZN(new_n1534));
  INV_X1    g1470(.A(new_n1534), .ZN(new_n1535));
  NOR2_X1   g1471(.A1(new_n1482), .A2(new_n1535), .ZN(new_n1536));
  AOI21_X1  g1472(.A(new_n1536), .B1(new_n1482), .B2(new_n1535), .ZN(new_n1537));
  INV_X1    g1473(.A(new_n1537), .ZN(new_n1538));
  NOR2_X1   g1474(.A1(new_n1452), .A2(new_n1455), .ZN(new_n1539));
  NOR2_X1   g1475(.A1(new_n1538), .A2(new_n1539), .ZN(new_n1540));
  AOI21_X1  g1476(.A(new_n1540), .B1(new_n1538), .B2(new_n1539), .ZN(new_n1541));
  INV_X1    g1477(.A(new_n1541), .ZN(new_n1542));
  NOR2_X1   g1478(.A1(new_n1481), .A2(new_n1542), .ZN(new_n1543));
  AOI21_X1  g1479(.A(new_n1543), .B1(new_n1481), .B2(new_n1542), .ZN(new_n1544));
  INV_X1    g1480(.A(new_n1544), .ZN(new_n1545));
  NOR2_X1   g1481(.A1(new_n1459), .A2(new_n1462), .ZN(new_n1546));
  NOR2_X1   g1482(.A1(new_n1545), .A2(new_n1546), .ZN(new_n1547));
  AOI21_X1  g1483(.A(new_n1547), .B1(new_n1545), .B2(new_n1546), .ZN(new_n1548));
  INV_X1    g1484(.A(new_n1548), .ZN(new_n1549));
  NOR2_X1   g1485(.A1(new_n1480), .A2(new_n1549), .ZN(new_n1550));
  AOI21_X1  g1486(.A(new_n1550), .B1(new_n1480), .B2(new_n1549), .ZN(new_n1551));
  INV_X1    g1487(.A(new_n1551), .ZN(new_n1552));
  NOR2_X1   g1488(.A1(new_n1466), .A2(new_n1469), .ZN(new_n1553));
  NOR2_X1   g1489(.A1(new_n1552), .A2(new_n1553), .ZN(new_n1554));
  AOI21_X1  g1490(.A(new_n1554), .B1(new_n1552), .B2(new_n1553), .ZN(new_n1555));
  INV_X1    g1491(.A(new_n1555), .ZN(new_n1556));
  NOR2_X1   g1492(.A1(new_n1479), .A2(new_n1556), .ZN(new_n1557));
  AOI21_X1  g1493(.A(new_n1557), .B1(new_n1479), .B2(new_n1556), .ZN(new_n1558));
  INV_X1    g1494(.A(new_n1558), .ZN(G6278));
  NOR2_X1   g1495(.A1(new_n1554), .A2(new_n1557), .ZN(new_n1560));
  NOR2_X1   g1496(.A1(new_n221), .A2(new_n854), .ZN(new_n1561));
  NOR2_X1   g1497(.A1(new_n274), .A2(new_n744), .ZN(new_n1562));
  NOR2_X1   g1498(.A1(new_n335), .A2(new_n644), .ZN(new_n1563));
  NOR2_X1   g1499(.A1(new_n404), .A2(new_n552), .ZN(new_n1564));
  NOR2_X1   g1500(.A1(new_n481), .A2(new_n468), .ZN(new_n1565));
  NOR2_X1   g1501(.A1(new_n566), .A2(new_n392), .ZN(new_n1566));
  NOR2_X1   g1502(.A1(new_n659), .A2(new_n324), .ZN(new_n1567));
  NOR2_X1   g1503(.A1(new_n760), .A2(new_n264), .ZN(new_n1568));
  NOR2_X1   g1504(.A1(new_n869), .A2(new_n212), .ZN(new_n1569));
  NOR2_X1   g1505(.A1(new_n1491), .A2(new_n1494), .ZN(new_n1570));
  NOR2_X1   g1506(.A1(new_n1569), .A2(new_n1570), .ZN(new_n1571));
  AOI21_X1  g1507(.A(new_n1571), .B1(new_n1569), .B2(new_n1570), .ZN(new_n1572));
  INV_X1    g1508(.A(new_n1572), .ZN(new_n1573));
  NOR2_X1   g1509(.A1(new_n1568), .A2(new_n1573), .ZN(new_n1574));
  AOI21_X1  g1510(.A(new_n1574), .B1(new_n1568), .B2(new_n1573), .ZN(new_n1575));
  INV_X1    g1511(.A(new_n1575), .ZN(new_n1576));
  NOR2_X1   g1512(.A1(new_n1498), .A2(new_n1501), .ZN(new_n1577));
  NOR2_X1   g1513(.A1(new_n1576), .A2(new_n1577), .ZN(new_n1578));
  AOI21_X1  g1514(.A(new_n1578), .B1(new_n1576), .B2(new_n1577), .ZN(new_n1579));
  INV_X1    g1515(.A(new_n1579), .ZN(new_n1580));
  NOR2_X1   g1516(.A1(new_n1567), .A2(new_n1580), .ZN(new_n1581));
  AOI21_X1  g1517(.A(new_n1581), .B1(new_n1567), .B2(new_n1580), .ZN(new_n1582));
  INV_X1    g1518(.A(new_n1582), .ZN(new_n1583));
  NOR2_X1   g1519(.A1(new_n1505), .A2(new_n1508), .ZN(new_n1584));
  NOR2_X1   g1520(.A1(new_n1583), .A2(new_n1584), .ZN(new_n1585));
  AOI21_X1  g1521(.A(new_n1585), .B1(new_n1583), .B2(new_n1584), .ZN(new_n1586));
  INV_X1    g1522(.A(new_n1586), .ZN(new_n1587));
  NOR2_X1   g1523(.A1(new_n1566), .A2(new_n1587), .ZN(new_n1588));
  AOI21_X1  g1524(.A(new_n1588), .B1(new_n1566), .B2(new_n1587), .ZN(new_n1589));
  INV_X1    g1525(.A(new_n1589), .ZN(new_n1590));
  NOR2_X1   g1526(.A1(new_n1512), .A2(new_n1515), .ZN(new_n1591));
  NOR2_X1   g1527(.A1(new_n1590), .A2(new_n1591), .ZN(new_n1592));
  AOI21_X1  g1528(.A(new_n1592), .B1(new_n1590), .B2(new_n1591), .ZN(new_n1593));
  INV_X1    g1529(.A(new_n1593), .ZN(new_n1594));
  NOR2_X1   g1530(.A1(new_n1565), .A2(new_n1594), .ZN(new_n1595));
  AOI21_X1  g1531(.A(new_n1595), .B1(new_n1565), .B2(new_n1594), .ZN(new_n1596));
  INV_X1    g1532(.A(new_n1596), .ZN(new_n1597));
  NOR2_X1   g1533(.A1(new_n1519), .A2(new_n1522), .ZN(new_n1598));
  NOR2_X1   g1534(.A1(new_n1597), .A2(new_n1598), .ZN(new_n1599));
  AOI21_X1  g1535(.A(new_n1599), .B1(new_n1597), .B2(new_n1598), .ZN(new_n1600));
  INV_X1    g1536(.A(new_n1600), .ZN(new_n1601));
  NOR2_X1   g1537(.A1(new_n1564), .A2(new_n1601), .ZN(new_n1602));
  AOI21_X1  g1538(.A(new_n1602), .B1(new_n1564), .B2(new_n1601), .ZN(new_n1603));
  INV_X1    g1539(.A(new_n1603), .ZN(new_n1604));
  NOR2_X1   g1540(.A1(new_n1526), .A2(new_n1529), .ZN(new_n1605));
  NOR2_X1   g1541(.A1(new_n1604), .A2(new_n1605), .ZN(new_n1606));
  AOI21_X1  g1542(.A(new_n1606), .B1(new_n1604), .B2(new_n1605), .ZN(new_n1607));
  INV_X1    g1543(.A(new_n1607), .ZN(new_n1608));
  NOR2_X1   g1544(.A1(new_n1563), .A2(new_n1608), .ZN(new_n1609));
  AOI21_X1  g1545(.A(new_n1609), .B1(new_n1563), .B2(new_n1608), .ZN(new_n1610));
  INV_X1    g1546(.A(new_n1610), .ZN(new_n1611));
  NOR2_X1   g1547(.A1(new_n1533), .A2(new_n1536), .ZN(new_n1612));
  NOR2_X1   g1548(.A1(new_n1611), .A2(new_n1612), .ZN(new_n1613));
  AOI21_X1  g1549(.A(new_n1613), .B1(new_n1611), .B2(new_n1612), .ZN(new_n1614));
  INV_X1    g1550(.A(new_n1614), .ZN(new_n1615));
  NOR2_X1   g1551(.A1(new_n1562), .A2(new_n1615), .ZN(new_n1616));
  AOI21_X1  g1552(.A(new_n1616), .B1(new_n1562), .B2(new_n1615), .ZN(new_n1617));
  INV_X1    g1553(.A(new_n1617), .ZN(new_n1618));
  NOR2_X1   g1554(.A1(new_n1540), .A2(new_n1543), .ZN(new_n1619));
  NOR2_X1   g1555(.A1(new_n1618), .A2(new_n1619), .ZN(new_n1620));
  AOI21_X1  g1556(.A(new_n1620), .B1(new_n1618), .B2(new_n1619), .ZN(new_n1621));
  INV_X1    g1557(.A(new_n1621), .ZN(new_n1622));
  NOR2_X1   g1558(.A1(new_n1561), .A2(new_n1622), .ZN(new_n1623));
  AOI21_X1  g1559(.A(new_n1623), .B1(new_n1561), .B2(new_n1622), .ZN(new_n1624));
  INV_X1    g1560(.A(new_n1624), .ZN(new_n1625));
  NOR2_X1   g1561(.A1(new_n1547), .A2(new_n1550), .ZN(new_n1626));
  NOR2_X1   g1562(.A1(new_n1625), .A2(new_n1626), .ZN(new_n1627));
  AOI21_X1  g1563(.A(new_n1627), .B1(new_n1625), .B2(new_n1626), .ZN(new_n1628));
  INV_X1    g1564(.A(new_n1628), .ZN(new_n1629));
  NOR2_X1   g1565(.A1(new_n1560), .A2(new_n1629), .ZN(new_n1630));
  AOI21_X1  g1566(.A(new_n1630), .B1(new_n1560), .B2(new_n1629), .ZN(new_n1631));
  INV_X1    g1567(.A(new_n1631), .ZN(G6279));
  NOR2_X1   g1568(.A1(new_n1627), .A2(new_n1630), .ZN(new_n1633));
  NOR2_X1   g1569(.A1(new_n274), .A2(new_n854), .ZN(new_n1634));
  NOR2_X1   g1570(.A1(new_n335), .A2(new_n744), .ZN(new_n1635));
  NOR2_X1   g1571(.A1(new_n404), .A2(new_n644), .ZN(new_n1636));
  NOR2_X1   g1572(.A1(new_n481), .A2(new_n552), .ZN(new_n1637));
  NOR2_X1   g1573(.A1(new_n566), .A2(new_n468), .ZN(new_n1638));
  NOR2_X1   g1574(.A1(new_n659), .A2(new_n392), .ZN(new_n1639));
  NOR2_X1   g1575(.A1(new_n760), .A2(new_n324), .ZN(new_n1640));
  NOR2_X1   g1576(.A1(new_n869), .A2(new_n264), .ZN(new_n1641));
  NOR2_X1   g1577(.A1(new_n1571), .A2(new_n1574), .ZN(new_n1642));
  NOR2_X1   g1578(.A1(new_n1641), .A2(new_n1642), .ZN(new_n1643));
  AOI21_X1  g1579(.A(new_n1643), .B1(new_n1641), .B2(new_n1642), .ZN(new_n1644));
  INV_X1    g1580(.A(new_n1644), .ZN(new_n1645));
  NOR2_X1   g1581(.A1(new_n1640), .A2(new_n1645), .ZN(new_n1646));
  AOI21_X1  g1582(.A(new_n1646), .B1(new_n1640), .B2(new_n1645), .ZN(new_n1647));
  INV_X1    g1583(.A(new_n1647), .ZN(new_n1648));
  NOR2_X1   g1584(.A1(new_n1578), .A2(new_n1581), .ZN(new_n1649));
  NOR2_X1   g1585(.A1(new_n1648), .A2(new_n1649), .ZN(new_n1650));
  AOI21_X1  g1586(.A(new_n1650), .B1(new_n1648), .B2(new_n1649), .ZN(new_n1651));
  INV_X1    g1587(.A(new_n1651), .ZN(new_n1652));
  NOR2_X1   g1588(.A1(new_n1639), .A2(new_n1652), .ZN(new_n1653));
  AOI21_X1  g1589(.A(new_n1653), .B1(new_n1639), .B2(new_n1652), .ZN(new_n1654));
  INV_X1    g1590(.A(new_n1654), .ZN(new_n1655));
  NOR2_X1   g1591(.A1(new_n1585), .A2(new_n1588), .ZN(new_n1656));
  NOR2_X1   g1592(.A1(new_n1655), .A2(new_n1656), .ZN(new_n1657));
  AOI21_X1  g1593(.A(new_n1657), .B1(new_n1655), .B2(new_n1656), .ZN(new_n1658));
  INV_X1    g1594(.A(new_n1658), .ZN(new_n1659));
  NOR2_X1   g1595(.A1(new_n1638), .A2(new_n1659), .ZN(new_n1660));
  AOI21_X1  g1596(.A(new_n1660), .B1(new_n1638), .B2(new_n1659), .ZN(new_n1661));
  INV_X1    g1597(.A(new_n1661), .ZN(new_n1662));
  NOR2_X1   g1598(.A1(new_n1592), .A2(new_n1595), .ZN(new_n1663));
  NOR2_X1   g1599(.A1(new_n1662), .A2(new_n1663), .ZN(new_n1664));
  AOI21_X1  g1600(.A(new_n1664), .B1(new_n1662), .B2(new_n1663), .ZN(new_n1665));
  INV_X1    g1601(.A(new_n1665), .ZN(new_n1666));
  NOR2_X1   g1602(.A1(new_n1637), .A2(new_n1666), .ZN(new_n1667));
  AOI21_X1  g1603(.A(new_n1667), .B1(new_n1637), .B2(new_n1666), .ZN(new_n1668));
  INV_X1    g1604(.A(new_n1668), .ZN(new_n1669));
  NOR2_X1   g1605(.A1(new_n1599), .A2(new_n1602), .ZN(new_n1670));
  NOR2_X1   g1606(.A1(new_n1669), .A2(new_n1670), .ZN(new_n1671));
  AOI21_X1  g1607(.A(new_n1671), .B1(new_n1669), .B2(new_n1670), .ZN(new_n1672));
  INV_X1    g1608(.A(new_n1672), .ZN(new_n1673));
  NOR2_X1   g1609(.A1(new_n1636), .A2(new_n1673), .ZN(new_n1674));
  AOI21_X1  g1610(.A(new_n1674), .B1(new_n1636), .B2(new_n1673), .ZN(new_n1675));
  INV_X1    g1611(.A(new_n1675), .ZN(new_n1676));
  NOR2_X1   g1612(.A1(new_n1606), .A2(new_n1609), .ZN(new_n1677));
  NOR2_X1   g1613(.A1(new_n1676), .A2(new_n1677), .ZN(new_n1678));
  AOI21_X1  g1614(.A(new_n1678), .B1(new_n1676), .B2(new_n1677), .ZN(new_n1679));
  INV_X1    g1615(.A(new_n1679), .ZN(new_n1680));
  NOR2_X1   g1616(.A1(new_n1635), .A2(new_n1680), .ZN(new_n1681));
  AOI21_X1  g1617(.A(new_n1681), .B1(new_n1635), .B2(new_n1680), .ZN(new_n1682));
  INV_X1    g1618(.A(new_n1682), .ZN(new_n1683));
  NOR2_X1   g1619(.A1(new_n1613), .A2(new_n1616), .ZN(new_n1684));
  NOR2_X1   g1620(.A1(new_n1683), .A2(new_n1684), .ZN(new_n1685));
  AOI21_X1  g1621(.A(new_n1685), .B1(new_n1683), .B2(new_n1684), .ZN(new_n1686));
  INV_X1    g1622(.A(new_n1686), .ZN(new_n1687));
  NOR2_X1   g1623(.A1(new_n1634), .A2(new_n1687), .ZN(new_n1688));
  AOI21_X1  g1624(.A(new_n1688), .B1(new_n1634), .B2(new_n1687), .ZN(new_n1689));
  INV_X1    g1625(.A(new_n1689), .ZN(new_n1690));
  NOR2_X1   g1626(.A1(new_n1620), .A2(new_n1623), .ZN(new_n1691));
  NOR2_X1   g1627(.A1(new_n1690), .A2(new_n1691), .ZN(new_n1692));
  AOI21_X1  g1628(.A(new_n1692), .B1(new_n1690), .B2(new_n1691), .ZN(new_n1693));
  INV_X1    g1629(.A(new_n1693), .ZN(new_n1694));
  NOR2_X1   g1630(.A1(new_n1633), .A2(new_n1694), .ZN(new_n1695));
  AOI21_X1  g1631(.A(new_n1695), .B1(new_n1633), .B2(new_n1694), .ZN(new_n1696));
  INV_X1    g1632(.A(new_n1696), .ZN(G6280));
  NOR2_X1   g1633(.A1(new_n1692), .A2(new_n1695), .ZN(new_n1698));
  NOR2_X1   g1634(.A1(new_n335), .A2(new_n854), .ZN(new_n1699));
  NOR2_X1   g1635(.A1(new_n404), .A2(new_n744), .ZN(new_n1700));
  NOR2_X1   g1636(.A1(new_n481), .A2(new_n644), .ZN(new_n1701));
  NOR2_X1   g1637(.A1(new_n566), .A2(new_n552), .ZN(new_n1702));
  NOR2_X1   g1638(.A1(new_n659), .A2(new_n468), .ZN(new_n1703));
  NOR2_X1   g1639(.A1(new_n760), .A2(new_n392), .ZN(new_n1704));
  NOR2_X1   g1640(.A1(new_n869), .A2(new_n324), .ZN(new_n1705));
  NOR2_X1   g1641(.A1(new_n1643), .A2(new_n1646), .ZN(new_n1706));
  NOR2_X1   g1642(.A1(new_n1705), .A2(new_n1706), .ZN(new_n1707));
  AOI21_X1  g1643(.A(new_n1707), .B1(new_n1705), .B2(new_n1706), .ZN(new_n1708));
  INV_X1    g1644(.A(new_n1708), .ZN(new_n1709));
  NOR2_X1   g1645(.A1(new_n1704), .A2(new_n1709), .ZN(new_n1710));
  AOI21_X1  g1646(.A(new_n1710), .B1(new_n1704), .B2(new_n1709), .ZN(new_n1711));
  INV_X1    g1647(.A(new_n1711), .ZN(new_n1712));
  NOR2_X1   g1648(.A1(new_n1650), .A2(new_n1653), .ZN(new_n1713));
  NOR2_X1   g1649(.A1(new_n1712), .A2(new_n1713), .ZN(new_n1714));
  AOI21_X1  g1650(.A(new_n1714), .B1(new_n1712), .B2(new_n1713), .ZN(new_n1715));
  INV_X1    g1651(.A(new_n1715), .ZN(new_n1716));
  NOR2_X1   g1652(.A1(new_n1703), .A2(new_n1716), .ZN(new_n1717));
  AOI21_X1  g1653(.A(new_n1717), .B1(new_n1703), .B2(new_n1716), .ZN(new_n1718));
  INV_X1    g1654(.A(new_n1718), .ZN(new_n1719));
  NOR2_X1   g1655(.A1(new_n1657), .A2(new_n1660), .ZN(new_n1720));
  NOR2_X1   g1656(.A1(new_n1719), .A2(new_n1720), .ZN(new_n1721));
  AOI21_X1  g1657(.A(new_n1721), .B1(new_n1719), .B2(new_n1720), .ZN(new_n1722));
  INV_X1    g1658(.A(new_n1722), .ZN(new_n1723));
  NOR2_X1   g1659(.A1(new_n1702), .A2(new_n1723), .ZN(new_n1724));
  AOI21_X1  g1660(.A(new_n1724), .B1(new_n1702), .B2(new_n1723), .ZN(new_n1725));
  INV_X1    g1661(.A(new_n1725), .ZN(new_n1726));
  NOR2_X1   g1662(.A1(new_n1664), .A2(new_n1667), .ZN(new_n1727));
  NOR2_X1   g1663(.A1(new_n1726), .A2(new_n1727), .ZN(new_n1728));
  AOI21_X1  g1664(.A(new_n1728), .B1(new_n1726), .B2(new_n1727), .ZN(new_n1729));
  INV_X1    g1665(.A(new_n1729), .ZN(new_n1730));
  NOR2_X1   g1666(.A1(new_n1701), .A2(new_n1730), .ZN(new_n1731));
  AOI21_X1  g1667(.A(new_n1731), .B1(new_n1701), .B2(new_n1730), .ZN(new_n1732));
  INV_X1    g1668(.A(new_n1732), .ZN(new_n1733));
  NOR2_X1   g1669(.A1(new_n1671), .A2(new_n1674), .ZN(new_n1734));
  NOR2_X1   g1670(.A1(new_n1733), .A2(new_n1734), .ZN(new_n1735));
  AOI21_X1  g1671(.A(new_n1735), .B1(new_n1733), .B2(new_n1734), .ZN(new_n1736));
  INV_X1    g1672(.A(new_n1736), .ZN(new_n1737));
  NOR2_X1   g1673(.A1(new_n1700), .A2(new_n1737), .ZN(new_n1738));
  AOI21_X1  g1674(.A(new_n1738), .B1(new_n1700), .B2(new_n1737), .ZN(new_n1739));
  INV_X1    g1675(.A(new_n1739), .ZN(new_n1740));
  NOR2_X1   g1676(.A1(new_n1678), .A2(new_n1681), .ZN(new_n1741));
  NOR2_X1   g1677(.A1(new_n1740), .A2(new_n1741), .ZN(new_n1742));
  AOI21_X1  g1678(.A(new_n1742), .B1(new_n1740), .B2(new_n1741), .ZN(new_n1743));
  INV_X1    g1679(.A(new_n1743), .ZN(new_n1744));
  NOR2_X1   g1680(.A1(new_n1699), .A2(new_n1744), .ZN(new_n1745));
  AOI21_X1  g1681(.A(new_n1745), .B1(new_n1699), .B2(new_n1744), .ZN(new_n1746));
  INV_X1    g1682(.A(new_n1746), .ZN(new_n1747));
  NOR2_X1   g1683(.A1(new_n1685), .A2(new_n1688), .ZN(new_n1748));
  NOR2_X1   g1684(.A1(new_n1747), .A2(new_n1748), .ZN(new_n1749));
  AOI21_X1  g1685(.A(new_n1749), .B1(new_n1747), .B2(new_n1748), .ZN(new_n1750));
  INV_X1    g1686(.A(new_n1750), .ZN(new_n1751));
  NOR2_X1   g1687(.A1(new_n1698), .A2(new_n1751), .ZN(new_n1752));
  AOI21_X1  g1688(.A(new_n1752), .B1(new_n1698), .B2(new_n1751), .ZN(new_n1753));
  INV_X1    g1689(.A(new_n1753), .ZN(G6281));
  NOR2_X1   g1690(.A1(new_n1749), .A2(new_n1752), .ZN(new_n1755));
  NOR2_X1   g1691(.A1(new_n404), .A2(new_n854), .ZN(new_n1756));
  NOR2_X1   g1692(.A1(new_n481), .A2(new_n744), .ZN(new_n1757));
  NOR2_X1   g1693(.A1(new_n566), .A2(new_n644), .ZN(new_n1758));
  NOR2_X1   g1694(.A1(new_n659), .A2(new_n552), .ZN(new_n1759));
  NOR2_X1   g1695(.A1(new_n760), .A2(new_n468), .ZN(new_n1760));
  NOR2_X1   g1696(.A1(new_n869), .A2(new_n392), .ZN(new_n1761));
  NOR2_X1   g1697(.A1(new_n1707), .A2(new_n1710), .ZN(new_n1762));
  NOR2_X1   g1698(.A1(new_n1761), .A2(new_n1762), .ZN(new_n1763));
  AOI21_X1  g1699(.A(new_n1763), .B1(new_n1761), .B2(new_n1762), .ZN(new_n1764));
  INV_X1    g1700(.A(new_n1764), .ZN(new_n1765));
  NOR2_X1   g1701(.A1(new_n1760), .A2(new_n1765), .ZN(new_n1766));
  AOI21_X1  g1702(.A(new_n1766), .B1(new_n1760), .B2(new_n1765), .ZN(new_n1767));
  INV_X1    g1703(.A(new_n1767), .ZN(new_n1768));
  NOR2_X1   g1704(.A1(new_n1714), .A2(new_n1717), .ZN(new_n1769));
  NOR2_X1   g1705(.A1(new_n1768), .A2(new_n1769), .ZN(new_n1770));
  AOI21_X1  g1706(.A(new_n1770), .B1(new_n1768), .B2(new_n1769), .ZN(new_n1771));
  INV_X1    g1707(.A(new_n1771), .ZN(new_n1772));
  NOR2_X1   g1708(.A1(new_n1759), .A2(new_n1772), .ZN(new_n1773));
  AOI21_X1  g1709(.A(new_n1773), .B1(new_n1759), .B2(new_n1772), .ZN(new_n1774));
  INV_X1    g1710(.A(new_n1774), .ZN(new_n1775));
  NOR2_X1   g1711(.A1(new_n1721), .A2(new_n1724), .ZN(new_n1776));
  NOR2_X1   g1712(.A1(new_n1775), .A2(new_n1776), .ZN(new_n1777));
  AOI21_X1  g1713(.A(new_n1777), .B1(new_n1775), .B2(new_n1776), .ZN(new_n1778));
  INV_X1    g1714(.A(new_n1778), .ZN(new_n1779));
  NOR2_X1   g1715(.A1(new_n1758), .A2(new_n1779), .ZN(new_n1780));
  AOI21_X1  g1716(.A(new_n1780), .B1(new_n1758), .B2(new_n1779), .ZN(new_n1781));
  INV_X1    g1717(.A(new_n1781), .ZN(new_n1782));
  NOR2_X1   g1718(.A1(new_n1728), .A2(new_n1731), .ZN(new_n1783));
  NOR2_X1   g1719(.A1(new_n1782), .A2(new_n1783), .ZN(new_n1784));
  AOI21_X1  g1720(.A(new_n1784), .B1(new_n1782), .B2(new_n1783), .ZN(new_n1785));
  INV_X1    g1721(.A(new_n1785), .ZN(new_n1786));
  NOR2_X1   g1722(.A1(new_n1757), .A2(new_n1786), .ZN(new_n1787));
  AOI21_X1  g1723(.A(new_n1787), .B1(new_n1757), .B2(new_n1786), .ZN(new_n1788));
  INV_X1    g1724(.A(new_n1788), .ZN(new_n1789));
  NOR2_X1   g1725(.A1(new_n1735), .A2(new_n1738), .ZN(new_n1790));
  NOR2_X1   g1726(.A1(new_n1789), .A2(new_n1790), .ZN(new_n1791));
  AOI21_X1  g1727(.A(new_n1791), .B1(new_n1789), .B2(new_n1790), .ZN(new_n1792));
  INV_X1    g1728(.A(new_n1792), .ZN(new_n1793));
  NOR2_X1   g1729(.A1(new_n1756), .A2(new_n1793), .ZN(new_n1794));
  AOI21_X1  g1730(.A(new_n1794), .B1(new_n1756), .B2(new_n1793), .ZN(new_n1795));
  INV_X1    g1731(.A(new_n1795), .ZN(new_n1796));
  NOR2_X1   g1732(.A1(new_n1742), .A2(new_n1745), .ZN(new_n1797));
  NOR2_X1   g1733(.A1(new_n1796), .A2(new_n1797), .ZN(new_n1798));
  AOI21_X1  g1734(.A(new_n1798), .B1(new_n1796), .B2(new_n1797), .ZN(new_n1799));
  INV_X1    g1735(.A(new_n1799), .ZN(new_n1800));
  NOR2_X1   g1736(.A1(new_n1755), .A2(new_n1800), .ZN(new_n1801));
  AOI21_X1  g1737(.A(new_n1801), .B1(new_n1755), .B2(new_n1800), .ZN(new_n1802));
  INV_X1    g1738(.A(new_n1802), .ZN(G6282));
  NOR2_X1   g1739(.A1(new_n1798), .A2(new_n1801), .ZN(new_n1804));
  NOR2_X1   g1740(.A1(new_n481), .A2(new_n854), .ZN(new_n1805));
  NOR2_X1   g1741(.A1(new_n566), .A2(new_n744), .ZN(new_n1806));
  NOR2_X1   g1742(.A1(new_n659), .A2(new_n644), .ZN(new_n1807));
  NOR2_X1   g1743(.A1(new_n760), .A2(new_n552), .ZN(new_n1808));
  NOR2_X1   g1744(.A1(new_n869), .A2(new_n468), .ZN(new_n1809));
  NOR2_X1   g1745(.A1(new_n1763), .A2(new_n1766), .ZN(new_n1810));
  NOR2_X1   g1746(.A1(new_n1809), .A2(new_n1810), .ZN(new_n1811));
  AOI21_X1  g1747(.A(new_n1811), .B1(new_n1809), .B2(new_n1810), .ZN(new_n1812));
  INV_X1    g1748(.A(new_n1812), .ZN(new_n1813));
  NOR2_X1   g1749(.A1(new_n1808), .A2(new_n1813), .ZN(new_n1814));
  AOI21_X1  g1750(.A(new_n1814), .B1(new_n1808), .B2(new_n1813), .ZN(new_n1815));
  INV_X1    g1751(.A(new_n1815), .ZN(new_n1816));
  NOR2_X1   g1752(.A1(new_n1770), .A2(new_n1773), .ZN(new_n1817));
  NOR2_X1   g1753(.A1(new_n1816), .A2(new_n1817), .ZN(new_n1818));
  AOI21_X1  g1754(.A(new_n1818), .B1(new_n1816), .B2(new_n1817), .ZN(new_n1819));
  INV_X1    g1755(.A(new_n1819), .ZN(new_n1820));
  NOR2_X1   g1756(.A1(new_n1807), .A2(new_n1820), .ZN(new_n1821));
  AOI21_X1  g1757(.A(new_n1821), .B1(new_n1807), .B2(new_n1820), .ZN(new_n1822));
  INV_X1    g1758(.A(new_n1822), .ZN(new_n1823));
  NOR2_X1   g1759(.A1(new_n1777), .A2(new_n1780), .ZN(new_n1824));
  NOR2_X1   g1760(.A1(new_n1823), .A2(new_n1824), .ZN(new_n1825));
  AOI21_X1  g1761(.A(new_n1825), .B1(new_n1823), .B2(new_n1824), .ZN(new_n1826));
  INV_X1    g1762(.A(new_n1826), .ZN(new_n1827));
  NOR2_X1   g1763(.A1(new_n1806), .A2(new_n1827), .ZN(new_n1828));
  AOI21_X1  g1764(.A(new_n1828), .B1(new_n1806), .B2(new_n1827), .ZN(new_n1829));
  INV_X1    g1765(.A(new_n1829), .ZN(new_n1830));
  NOR2_X1   g1766(.A1(new_n1784), .A2(new_n1787), .ZN(new_n1831));
  NOR2_X1   g1767(.A1(new_n1830), .A2(new_n1831), .ZN(new_n1832));
  AOI21_X1  g1768(.A(new_n1832), .B1(new_n1830), .B2(new_n1831), .ZN(new_n1833));
  INV_X1    g1769(.A(new_n1833), .ZN(new_n1834));
  NOR2_X1   g1770(.A1(new_n1805), .A2(new_n1834), .ZN(new_n1835));
  AOI21_X1  g1771(.A(new_n1835), .B1(new_n1805), .B2(new_n1834), .ZN(new_n1836));
  INV_X1    g1772(.A(new_n1836), .ZN(new_n1837));
  NOR2_X1   g1773(.A1(new_n1791), .A2(new_n1794), .ZN(new_n1838));
  NOR2_X1   g1774(.A1(new_n1837), .A2(new_n1838), .ZN(new_n1839));
  AOI21_X1  g1775(.A(new_n1839), .B1(new_n1837), .B2(new_n1838), .ZN(new_n1840));
  INV_X1    g1776(.A(new_n1840), .ZN(new_n1841));
  NOR2_X1   g1777(.A1(new_n1804), .A2(new_n1841), .ZN(new_n1842));
  AOI21_X1  g1778(.A(new_n1842), .B1(new_n1804), .B2(new_n1841), .ZN(new_n1843));
  INV_X1    g1779(.A(new_n1843), .ZN(G6283));
  NOR2_X1   g1780(.A1(new_n1839), .A2(new_n1842), .ZN(new_n1845));
  NOR2_X1   g1781(.A1(new_n566), .A2(new_n854), .ZN(new_n1846));
  NOR2_X1   g1782(.A1(new_n659), .A2(new_n744), .ZN(new_n1847));
  NOR2_X1   g1783(.A1(new_n760), .A2(new_n644), .ZN(new_n1848));
  NOR2_X1   g1784(.A1(new_n869), .A2(new_n552), .ZN(new_n1849));
  NOR2_X1   g1785(.A1(new_n1811), .A2(new_n1814), .ZN(new_n1850));
  NOR2_X1   g1786(.A1(new_n1849), .A2(new_n1850), .ZN(new_n1851));
  AOI21_X1  g1787(.A(new_n1851), .B1(new_n1849), .B2(new_n1850), .ZN(new_n1852));
  INV_X1    g1788(.A(new_n1852), .ZN(new_n1853));
  NOR2_X1   g1789(.A1(new_n1848), .A2(new_n1853), .ZN(new_n1854));
  AOI21_X1  g1790(.A(new_n1854), .B1(new_n1848), .B2(new_n1853), .ZN(new_n1855));
  INV_X1    g1791(.A(new_n1855), .ZN(new_n1856));
  NOR2_X1   g1792(.A1(new_n1818), .A2(new_n1821), .ZN(new_n1857));
  NOR2_X1   g1793(.A1(new_n1856), .A2(new_n1857), .ZN(new_n1858));
  AOI21_X1  g1794(.A(new_n1858), .B1(new_n1856), .B2(new_n1857), .ZN(new_n1859));
  INV_X1    g1795(.A(new_n1859), .ZN(new_n1860));
  NOR2_X1   g1796(.A1(new_n1847), .A2(new_n1860), .ZN(new_n1861));
  AOI21_X1  g1797(.A(new_n1861), .B1(new_n1847), .B2(new_n1860), .ZN(new_n1862));
  INV_X1    g1798(.A(new_n1862), .ZN(new_n1863));
  NOR2_X1   g1799(.A1(new_n1825), .A2(new_n1828), .ZN(new_n1864));
  NOR2_X1   g1800(.A1(new_n1863), .A2(new_n1864), .ZN(new_n1865));
  AOI21_X1  g1801(.A(new_n1865), .B1(new_n1863), .B2(new_n1864), .ZN(new_n1866));
  INV_X1    g1802(.A(new_n1866), .ZN(new_n1867));
  NOR2_X1   g1803(.A1(new_n1846), .A2(new_n1867), .ZN(new_n1868));
  AOI21_X1  g1804(.A(new_n1868), .B1(new_n1846), .B2(new_n1867), .ZN(new_n1869));
  INV_X1    g1805(.A(new_n1869), .ZN(new_n1870));
  NOR2_X1   g1806(.A1(new_n1832), .A2(new_n1835), .ZN(new_n1871));
  NOR2_X1   g1807(.A1(new_n1870), .A2(new_n1871), .ZN(new_n1872));
  AOI21_X1  g1808(.A(new_n1872), .B1(new_n1870), .B2(new_n1871), .ZN(new_n1873));
  INV_X1    g1809(.A(new_n1873), .ZN(new_n1874));
  NOR2_X1   g1810(.A1(new_n1845), .A2(new_n1874), .ZN(new_n1875));
  AOI21_X1  g1811(.A(new_n1875), .B1(new_n1845), .B2(new_n1874), .ZN(new_n1876));
  INV_X1    g1812(.A(new_n1876), .ZN(G6284));
  NOR2_X1   g1813(.A1(new_n1872), .A2(new_n1875), .ZN(new_n1878));
  NOR2_X1   g1814(.A1(new_n659), .A2(new_n854), .ZN(new_n1879));
  NOR2_X1   g1815(.A1(new_n760), .A2(new_n744), .ZN(new_n1880));
  NOR2_X1   g1816(.A1(new_n869), .A2(new_n644), .ZN(new_n1881));
  NOR2_X1   g1817(.A1(new_n1851), .A2(new_n1854), .ZN(new_n1882));
  NOR2_X1   g1818(.A1(new_n1881), .A2(new_n1882), .ZN(new_n1883));
  AOI21_X1  g1819(.A(new_n1883), .B1(new_n1881), .B2(new_n1882), .ZN(new_n1884));
  INV_X1    g1820(.A(new_n1884), .ZN(new_n1885));
  NOR2_X1   g1821(.A1(new_n1880), .A2(new_n1885), .ZN(new_n1886));
  AOI21_X1  g1822(.A(new_n1886), .B1(new_n1880), .B2(new_n1885), .ZN(new_n1887));
  INV_X1    g1823(.A(new_n1887), .ZN(new_n1888));
  NOR2_X1   g1824(.A1(new_n1858), .A2(new_n1861), .ZN(new_n1889));
  NOR2_X1   g1825(.A1(new_n1888), .A2(new_n1889), .ZN(new_n1890));
  AOI21_X1  g1826(.A(new_n1890), .B1(new_n1888), .B2(new_n1889), .ZN(new_n1891));
  INV_X1    g1827(.A(new_n1891), .ZN(new_n1892));
  NOR2_X1   g1828(.A1(new_n1879), .A2(new_n1892), .ZN(new_n1893));
  AOI21_X1  g1829(.A(new_n1893), .B1(new_n1879), .B2(new_n1892), .ZN(new_n1894));
  INV_X1    g1830(.A(new_n1894), .ZN(new_n1895));
  NOR2_X1   g1831(.A1(new_n1865), .A2(new_n1868), .ZN(new_n1896));
  NOR2_X1   g1832(.A1(new_n1895), .A2(new_n1896), .ZN(new_n1897));
  AOI21_X1  g1833(.A(new_n1897), .B1(new_n1895), .B2(new_n1896), .ZN(new_n1898));
  INV_X1    g1834(.A(new_n1898), .ZN(new_n1899));
  NOR2_X1   g1835(.A1(new_n1878), .A2(new_n1899), .ZN(new_n1900));
  AOI21_X1  g1836(.A(new_n1900), .B1(new_n1878), .B2(new_n1899), .ZN(new_n1901));
  INV_X1    g1837(.A(new_n1901), .ZN(G6285));
  NOR2_X1   g1838(.A1(new_n1897), .A2(new_n1900), .ZN(new_n1903));
  NOR2_X1   g1839(.A1(new_n760), .A2(new_n854), .ZN(new_n1904));
  NOR2_X1   g1840(.A1(new_n869), .A2(new_n744), .ZN(new_n1905));
  NOR2_X1   g1841(.A1(new_n1883), .A2(new_n1886), .ZN(new_n1906));
  NOR2_X1   g1842(.A1(new_n1905), .A2(new_n1906), .ZN(new_n1907));
  AOI21_X1  g1843(.A(new_n1907), .B1(new_n1905), .B2(new_n1906), .ZN(new_n1908));
  INV_X1    g1844(.A(new_n1908), .ZN(new_n1909));
  NOR2_X1   g1845(.A1(new_n1904), .A2(new_n1909), .ZN(new_n1910));
  AOI21_X1  g1846(.A(new_n1910), .B1(new_n1904), .B2(new_n1909), .ZN(new_n1911));
  INV_X1    g1847(.A(new_n1911), .ZN(new_n1912));
  NOR2_X1   g1848(.A1(new_n1890), .A2(new_n1893), .ZN(new_n1913));
  NOR2_X1   g1849(.A1(new_n1912), .A2(new_n1913), .ZN(new_n1914));
  AOI21_X1  g1850(.A(new_n1914), .B1(new_n1912), .B2(new_n1913), .ZN(new_n1915));
  INV_X1    g1851(.A(new_n1915), .ZN(new_n1916));
  NOR2_X1   g1852(.A1(new_n1903), .A2(new_n1916), .ZN(new_n1917));
  AOI21_X1  g1853(.A(new_n1917), .B1(new_n1903), .B2(new_n1916), .ZN(new_n1918));
  INV_X1    g1854(.A(new_n1918), .ZN(G6286));
  NOR2_X1   g1855(.A1(new_n869), .A2(new_n854), .ZN(new_n1920));
  NOR2_X1   g1856(.A1(new_n1907), .A2(new_n1910), .ZN(new_n1921));
  NOR2_X1   g1857(.A1(new_n1920), .A2(new_n1921), .ZN(new_n1922));
  OR2_X1    g1858(.A1(new_n1914), .A2(new_n1917), .ZN(new_n1923));
  AOI21_X1  g1859(.A(new_n1922), .B1(new_n1920), .B2(new_n1921), .ZN(new_n1924));
  AOI21_X1  g1860(.A(new_n1922), .B1(new_n1923), .B2(new_n1924), .ZN(G6287));
  XNOR2_X1  g1861(.A(new_n1923), .B(new_n1924), .ZN(G6288));
endmodule


