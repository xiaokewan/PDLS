// Benchmark "iscas85-original/c5315" written by ABC on Sat Nov 18 15:15:55 2023

module c5315  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160,
    G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172,
    G173, G174, G175, G176, G177, G178,
    G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178;
  output G5193, G5194, G5195, G5196, G5197, G5198, G5199, G5200, G5201, G5202,
    G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212,
    G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222,
    G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232,
    G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242,
    G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252,
    G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262,
    G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272,
    G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282,
    G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292,
    G5293, G5294, G5295, G5296, G5297, G5298, G5299, G5300, G5301, G5302,
    G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312,
    G5313, G5314, G5315;
  wire new_n321, new_n331, new_n339, new_n344, new_n346, new_n348, new_n350,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n510, new_n511, new_n512, new_n513, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n712,
    new_n714, new_n716, new_n718, new_n720, new_n722, new_n724, new_n726,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n735, new_n736,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n757,
    new_n758, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n779, new_n780, new_n782, new_n783, new_n785, new_n787, new_n789,
    new_n791, new_n793, new_n795, new_n797, new_n799, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n819, new_n820, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n931, new_n933,
    new_n934, new_n936, new_n937;
  INV_X1    g000(.A(G66), .ZN(G5193));
  INV_X1    g001(.A(G113), .ZN(G5194));
  INV_X1    g002(.A(G165), .ZN(G5195));
  INV_X1    g003(.A(G151), .ZN(G5196));
  INV_X1    g004(.A(G127), .ZN(G5197));
  INV_X1    g005(.A(G131), .ZN(G5198));
  INV_X1    g006(.A(G153), .ZN(G5207));
  INV_X1    g007(.A(G156), .ZN(G5208));
  NOR2_X1   g008(.A1(G5207), .A2(G5208), .ZN(G5199));
  INV_X1    g009(.A(G152), .ZN(G5200));
  BUF_X1    g010(.A(G5196), .Z(G5201));
  BUF_X1    g011(.A(G5196), .Z(G5202));
  INV_X1    g012(.A(G125), .ZN(G5203));
  INV_X1    g013(.A(G129), .ZN(G5204));
  AND2_X1   g014(.A1(G66), .A2(G67), .ZN(G5205));
  INV_X1    g015(.A(G99), .ZN(G5206));
  INV_X1    g016(.A(G155), .ZN(G5209));
  AND2_X1   g017(.A1(G1), .A2(G134), .ZN(G5210));
  AND2_X1   g018(.A1(G63), .A2(G5195), .ZN(G5211));
  INV_X1    g019(.A(G164), .ZN(new_n321));
  NAND2_X1  g020(.A1(G11), .A2(new_n321), .ZN(G5212));
  NAND2_X1  g021(.A1(G136), .A2(G154), .ZN(G5213));
  BUF_X1    g022(.A(G64), .Z(G5214));
  BUF_X1    g023(.A(G66), .Z(G5215));
  BUF_X1    g024(.A(G1), .Z(G5216));
  BUF_X1    g025(.A(G152), .Z(G5217));
  BUF_X1    g026(.A(G114), .Z(G5218));
  BUF_X1    g027(.A(G152), .Z(G5219));
  NAND2_X1  g028(.A1(G11), .A2(G12), .ZN(G5221));
  INV_X1    g029(.A(G5221), .ZN(new_n331));
  NAND2_X1  g030(.A1(G65), .A2(new_n331), .ZN(G5220));
  INV_X1    g031(.A(G1), .ZN(G5222));
  BUF_X1    g032(.A(G5222), .Z(G5223));
  BUF_X1    g033(.A(G5222), .Z(G5224));
  BUF_X1    g034(.A(G5222), .Z(G5225));
  INV_X1    g035(.A(G114), .ZN(G5226));
  BUF_X1    g036(.A(G5226), .Z(G5227));
  INV_X1    g037(.A(G163), .ZN(new_n339));
  OAI221_X1 g038(.A(new_n331), .B1(G33), .B2(G163), .C1(G34), .C2(new_n339), .ZN(G5228));
  OAI221_X1 g039(.A(new_n331), .B1(G35), .B2(G163), .C1(G13), .C2(new_n339), .ZN(G5229));
  BUF_X1    g040(.A(G5229), .Z(G5230));
  NAND2_X1  g041(.A1(G32), .A2(new_n331), .ZN(G5231));
  AOI221_X1 g042(.A(G5221), .B1(G9), .B2(new_n339), .C1(G8), .C2(G163), .ZN(new_n344));
  NOR2_X1   g043(.A1(G5193), .A2(new_n344), .ZN(G5232));
  AOI221_X1 g044(.A(G5221), .B1(G30), .B2(new_n339), .C1(G10), .C2(G163), .ZN(new_n346));
  NOR2_X1   g045(.A1(G5193), .A2(new_n346), .ZN(G5233));
  AOI221_X1 g046(.A(G5221), .B1(G7), .B2(new_n339), .C1(G28), .C2(G163), .ZN(new_n348));
  NOR2_X1   g047(.A1(G5193), .A2(new_n348), .ZN(G5234));
  AOI221_X1 g048(.A(G5221), .B1(G29), .B2(new_n339), .C1(G31), .C2(G163), .ZN(new_n350));
  NOR2_X1   g049(.A1(G5193), .A2(new_n350), .ZN(G5235));
  INV_X1    g050(.A(G121), .ZN(new_n352));
  OAI221_X1 g051(.A(G147), .B1(G121), .B2(G169), .C1(new_n352), .C2(G168), .ZN(new_n353));
  INV_X1    g052(.A(G167), .ZN(new_n354));
  NOR2_X1   g053(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g054(.A(G147), .ZN(new_n356));
  INV_X1    g055(.A(G166), .ZN(new_n357));
  OAI21_X1  g056(.A(new_n356), .B1(G121), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g057(.A(new_n353), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g058(.A(G126), .ZN(new_n360));
  OAI221_X1 g059(.A(G149), .B1(G126), .B2(G169), .C1(new_n360), .C2(G168), .ZN(new_n361));
  NOR2_X1   g060(.A1(new_n360), .A2(new_n354), .ZN(new_n362));
  INV_X1    g061(.A(G149), .ZN(new_n363));
  OAI21_X1  g062(.A(new_n363), .B1(G126), .B2(new_n357), .ZN(new_n364));
  OAI21_X1  g063(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g064(.A(G101), .ZN(new_n366));
  INV_X1    g065(.A(G130), .ZN(new_n367));
  INV_X1    g066(.A(G100), .ZN(new_n368));
  OAI22_X1  g067(.A1(new_n366), .A2(new_n367), .B1(new_n368), .B2(G130), .ZN(new_n369));
  INV_X1    g068(.A(G148), .ZN(new_n370));
  INV_X1    g069(.A(G169), .ZN(new_n371));
  OAI22_X1  g070(.A1(G148), .A2(G166), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g071(.A(G115), .ZN(new_n373));
  OAI22_X1  g072(.A1(new_n366), .A2(new_n373), .B1(new_n368), .B2(G115), .ZN(new_n374));
  INV_X1    g073(.A(new_n374), .ZN(new_n375));
  INV_X1    g074(.A(G102), .ZN(new_n376));
  INV_X1    g075(.A(G98), .ZN(new_n377));
  OAI22_X1  g076(.A1(new_n376), .A2(G5194), .B1(new_n377), .B2(G113), .ZN(new_n378));
  NAND2_X1  g077(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g078(.A(G128), .ZN(new_n380));
  OAI221_X1 g079(.A(G150), .B1(G128), .B2(G169), .C1(new_n380), .C2(G168), .ZN(new_n381));
  NOR2_X1   g080(.A1(new_n380), .A2(new_n354), .ZN(new_n382));
  INV_X1    g081(.A(G150), .ZN(new_n383));
  OAI21_X1  g082(.A(new_n383), .B1(G128), .B2(new_n357), .ZN(new_n384));
  OAI21_X1  g083(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OR4_X1    g084(.A1(new_n369), .A2(new_n372), .A3(new_n379), .A4(new_n385), .ZN(new_n386));
  INV_X1    g085(.A(G146), .ZN(new_n387));
  INV_X1    g086(.A(G119), .ZN(new_n388));
  AOI221_X1 g087(.A(new_n387), .B1(new_n368), .B2(new_n388), .C1(new_n366), .C2(G119), .ZN(new_n389));
  AOI221_X1 g088(.A(G146), .B1(G98), .B2(new_n388), .C1(G102), .C2(G119), .ZN(new_n390));
  OR2_X1    g089(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g090(.A(G145), .ZN(new_n392));
  INV_X1    g091(.A(G117), .ZN(new_n393));
  AOI221_X1 g092(.A(new_n392), .B1(new_n368), .B2(new_n393), .C1(new_n366), .C2(G117), .ZN(new_n394));
  AOI221_X1 g093(.A(G145), .B1(G98), .B2(new_n393), .C1(G102), .C2(G117), .ZN(new_n395));
  OR2_X1    g094(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g095(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NOR4_X1   g096(.A1(new_n359), .A2(new_n365), .A3(new_n386), .A4(new_n397), .ZN(G5236));
  INV_X1    g097(.A(G105), .ZN(new_n399));
  OAI221_X1 g098(.A(G138), .B1(G105), .B2(G169), .C1(new_n399), .C2(G168), .ZN(new_n400));
  NOR2_X1   g099(.A1(new_n399), .A2(new_n354), .ZN(new_n401));
  INV_X1    g100(.A(G138), .ZN(new_n402));
  OAI21_X1  g101(.A(new_n402), .B1(G105), .B2(new_n357), .ZN(new_n403));
  OAI21_X1  g102(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g103(.A(G103), .ZN(new_n405));
  OAI221_X1 g104(.A(G137), .B1(G103), .B2(G169), .C1(new_n405), .C2(G168), .ZN(new_n406));
  NOR2_X1   g105(.A1(new_n405), .A2(new_n354), .ZN(new_n407));
  INV_X1    g106(.A(G137), .ZN(new_n408));
  OAI21_X1  g107(.A(new_n408), .B1(G103), .B2(new_n357), .ZN(new_n409));
  OAI21_X1  g108(.A(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g109(.A(G141), .ZN(new_n411));
  INV_X1    g110(.A(G96), .ZN(new_n412));
  OAI221_X1 g111(.A(new_n411), .B1(G96), .B2(G166), .C1(new_n412), .C2(G167), .ZN(new_n413));
  NAND2_X1  g112(.A1(new_n412), .A2(G141), .ZN(new_n414));
  NAND2_X1  g113(.A1(G96), .A2(G141), .ZN(new_n415));
  OAI221_X1 g114(.A(new_n413), .B1(G169), .B2(new_n414), .C1(G168), .C2(new_n415), .ZN(new_n416));
  INV_X1    g115(.A(new_n416), .ZN(new_n417));
  INV_X1    g116(.A(G109), .ZN(new_n418));
  OAI221_X1 g117(.A(G135), .B1(G109), .B2(G169), .C1(new_n418), .C2(G168), .ZN(new_n419));
  NOR2_X1   g118(.A1(new_n418), .A2(new_n354), .ZN(new_n420));
  INV_X1    g119(.A(G135), .ZN(new_n421));
  OAI21_X1  g120(.A(new_n421), .B1(G109), .B2(new_n357), .ZN(new_n422));
  OAI21_X1  g121(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g122(.A(G143), .ZN(new_n424));
  INV_X1    g123(.A(G90), .ZN(new_n425));
  OAI221_X1 g124(.A(new_n424), .B1(G90), .B2(G166), .C1(new_n425), .C2(G167), .ZN(new_n426));
  NAND2_X1  g125(.A1(new_n425), .A2(G143), .ZN(new_n427));
  NAND2_X1  g126(.A1(G90), .A2(G143), .ZN(new_n428));
  OAI221_X1 g127(.A(new_n426), .B1(G169), .B2(new_n427), .C1(G168), .C2(new_n428), .ZN(new_n429));
  INV_X1    g128(.A(new_n429), .ZN(new_n430));
  INV_X1    g129(.A(G107), .ZN(new_n431));
  OAI221_X1 g130(.A(G139), .B1(G107), .B2(G169), .C1(new_n431), .C2(G168), .ZN(new_n432));
  NOR2_X1   g131(.A1(new_n431), .A2(new_n354), .ZN(new_n433));
  INV_X1    g132(.A(G139), .ZN(new_n434));
  OAI21_X1  g133(.A(new_n434), .B1(G107), .B2(new_n357), .ZN(new_n435));
  OAI21_X1  g134(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g135(.A(new_n436), .ZN(new_n437));
  INV_X1    g136(.A(G140), .ZN(new_n438));
  INV_X1    g137(.A(G94), .ZN(new_n439));
  OAI221_X1 g138(.A(new_n438), .B1(G94), .B2(G166), .C1(new_n439), .C2(G167), .ZN(new_n440));
  NAND2_X1  g139(.A1(new_n439), .A2(G140), .ZN(new_n441));
  NAND2_X1  g140(.A1(G94), .A2(G140), .ZN(new_n442));
  OAI221_X1 g141(.A(new_n440), .B1(G169), .B2(new_n441), .C1(G168), .C2(new_n442), .ZN(new_n443));
  INV_X1    g142(.A(G142), .ZN(new_n444));
  INV_X1    g143(.A(G88), .ZN(new_n445));
  AOI221_X1 g144(.A(new_n444), .B1(new_n445), .B2(new_n366), .C1(G88), .C2(new_n368), .ZN(new_n446));
  AOI221_X1 g145(.A(G142), .B1(new_n445), .B2(G102), .C1(G88), .C2(G98), .ZN(new_n447));
  NOR2_X1   g146(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g147(.A(G144), .ZN(new_n449));
  INV_X1    g148(.A(G92), .ZN(new_n450));
  OAI221_X1 g149(.A(new_n449), .B1(G92), .B2(G166), .C1(new_n450), .C2(G167), .ZN(new_n451));
  NAND2_X1  g150(.A1(new_n450), .A2(G144), .ZN(new_n452));
  NAND2_X1  g151(.A1(G92), .A2(G144), .ZN(new_n453));
  OAI221_X1 g152(.A(new_n451), .B1(G169), .B2(new_n452), .C1(G168), .C2(new_n453), .ZN(new_n454));
  NAND4_X1  g153(.A1(new_n437), .A2(new_n443), .A3(new_n448), .A4(new_n454), .ZN(new_n455));
  OR3_X1    g154(.A1(new_n423), .A2(new_n430), .A3(new_n455), .ZN(new_n456));
  NOR4_X1   g155(.A1(new_n404), .A2(new_n410), .A3(new_n417), .A4(new_n456), .ZN(G5237));
  INV_X1    g156(.A(G124), .ZN(new_n458));
  OAI22_X1  g157(.A1(G104), .A2(G124), .B1(G103), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g158(.A1(new_n408), .A2(new_n459), .ZN(new_n460));
  INV_X1    g159(.A(new_n459), .ZN(new_n461));
  NOR2_X1   g160(.A1(G137), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g161(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g162(.A(new_n463), .ZN(new_n464));
  OAI22_X1  g163(.A1(G106), .A2(G124), .B1(G105), .B2(new_n458), .ZN(new_n465));
  NOR2_X1   g164(.A1(new_n402), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g165(.A1(new_n402), .A2(new_n465), .ZN(new_n467));
  NOR2_X1   g166(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g167(.A(new_n468), .ZN(new_n469));
  OAI22_X1  g168(.A1(G97), .A2(G124), .B1(G96), .B2(new_n458), .ZN(new_n470));
  NAND2_X1  g169(.A1(new_n411), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g170(.A(new_n471), .B1(new_n411), .B2(new_n470), .ZN(new_n472));
  OAI22_X1  g171(.A1(G108), .A2(G124), .B1(G107), .B2(new_n458), .ZN(new_n473));
  XNOR2_X1  g172(.A(new_n434), .B(new_n473), .ZN(new_n474));
  OAI22_X1  g173(.A1(G110), .A2(G124), .B1(G109), .B2(new_n458), .ZN(new_n475));
  NOR2_X1   g174(.A1(new_n421), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g175(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g176(.A(new_n475), .ZN(new_n478));
  OAI21_X1  g177(.A(new_n477), .B1(G135), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g178(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  OR3_X1    g179(.A1(new_n464), .A2(new_n469), .A3(new_n480), .ZN(new_n481));
  OAI22_X1  g180(.A1(G93), .A2(G124), .B1(G92), .B2(new_n458), .ZN(new_n482));
  OAI22_X1  g181(.A1(G95), .A2(G124), .B1(G94), .B2(new_n458), .ZN(new_n483));
  OR2_X1    g182(.A1(new_n438), .A2(new_n483), .ZN(new_n484));
  INV_X1    g183(.A(new_n482), .ZN(new_n485));
  OAI22_X1  g184(.A1(new_n449), .A2(new_n482), .B1(G144), .B2(new_n485), .ZN(new_n486));
  OAI22_X1  g185(.A1(new_n449), .A2(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g186(.A(new_n487), .ZN(new_n488));
  OAI22_X1  g187(.A1(G91), .A2(G124), .B1(G90), .B2(new_n458), .ZN(new_n489));
  INV_X1    g188(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g189(.A1(G143), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g190(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g191(.A1(new_n424), .A2(new_n489), .ZN(new_n493));
  INV_X1    g192(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g193(.A(new_n492), .B1(new_n494), .B2(new_n488), .ZN(new_n495));
  OAI22_X1  g194(.A1(G89), .A2(G124), .B1(G88), .B2(new_n458), .ZN(new_n496));
  INV_X1    g195(.A(new_n496), .ZN(new_n497));
  OAI22_X1  g196(.A1(new_n444), .A2(new_n496), .B1(G142), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g197(.A1(new_n438), .A2(new_n483), .ZN(new_n499));
  NAND2_X1  g198(.A1(new_n484), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g199(.A1(new_n486), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g200(.A(new_n484), .B(new_n486), .Z(new_n502));
  INV_X1    g201(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g202(.A(new_n501), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g203(.A(new_n498), .B(new_n504), .Z(new_n505));
  INV_X1    g204(.A(new_n491), .ZN(new_n506));
  NAND2_X1  g205(.A1(new_n506), .A2(new_n501), .ZN(new_n507));
  OR3_X1    g206(.A1(new_n495), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g207(.A1(new_n481), .A2(new_n508), .ZN(G5238));
  INV_X1    g208(.A(G123), .ZN(new_n510));
  OAI22_X1  g209(.A1(G114), .A2(G123), .B1(G113), .B2(new_n510), .ZN(new_n511));
  OAI22_X1  g210(.A1(G116), .A2(G123), .B1(G115), .B2(new_n510), .ZN(new_n512));
  INV_X1    g211(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g212(.A1(new_n511), .A2(new_n513), .ZN(G5245));
  OAI21_X1  g213(.A(G5245), .B1(new_n511), .B2(new_n513), .ZN(G5251));
  OAI22_X1  g214(.A1(G120), .A2(G123), .B1(G119), .B2(new_n510), .ZN(new_n516));
  INV_X1    g215(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g216(.A1(G146), .A2(new_n517), .ZN(new_n518));
  OAI22_X1  g217(.A1(G118), .A2(G123), .B1(G117), .B2(new_n510), .ZN(new_n519));
  AND2_X1   g218(.A1(new_n392), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g219(.A1(new_n387), .A2(new_n516), .ZN(new_n521));
  NOR2_X1   g220(.A1(new_n392), .A2(new_n519), .ZN(new_n522));
  INV_X1    g221(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g222(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g223(.A(new_n512), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g224(.A(new_n518), .B(new_n525), .ZN(new_n526));
  OAI22_X1  g225(.A1(G123), .A2(G127), .B1(new_n510), .B2(G126), .ZN(new_n527));
  NOR2_X1   g226(.A1(new_n363), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g227(.A1(new_n363), .A2(new_n527), .ZN(new_n529));
  OR2_X1    g228(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI22_X1  g229(.A1(G123), .A2(G129), .B1(new_n510), .B2(G128), .ZN(new_n531));
  NOR2_X1   g230(.A1(new_n383), .A2(new_n531), .ZN(new_n532));
  INV_X1    g231(.A(new_n532), .ZN(new_n533));
  OAI22_X1  g232(.A1(G123), .A2(G131), .B1(new_n510), .B2(G130), .ZN(new_n534));
  INV_X1    g233(.A(new_n531), .ZN(new_n535));
  OAI21_X1  g234(.A(new_n534), .B1(G150), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g235(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  OAI22_X1  g236(.A1(new_n363), .A2(new_n527), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g237(.A1(G123), .A2(G125), .ZN(new_n539));
  NOR2_X1   g238(.A1(new_n370), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g239(.A(new_n540), .B1(new_n370), .B2(new_n539), .ZN(new_n541));
  NAND2_X1  g240(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  OAI22_X1  g241(.A1(G122), .A2(G123), .B1(G121), .B2(new_n510), .ZN(new_n543));
  XOR2_X1   g242(.A(new_n356), .B(new_n543), .Z(new_n544));
  NOR2_X1   g243(.A1(new_n520), .A2(new_n522), .ZN(new_n545));
  OAI211_X1 g244(.A(new_n544), .B(new_n545), .C1(new_n529), .C2(new_n533), .ZN(new_n546));
  OR4_X1    g245(.A1(new_n518), .A2(new_n521), .A3(new_n528), .A4(new_n546), .ZN(new_n547));
  NOR4_X1   g246(.A1(G5251), .A2(new_n526), .A3(new_n542), .A4(new_n547), .ZN(G5239));
  BUF_X1    g247(.A(G5239), .Z(G5240));
  BUF_X1    g248(.A(G5238), .Z(G5241));
  OAI22_X1  g249(.A1(G126), .A2(G128), .B1(new_n360), .B2(new_n380), .ZN(new_n551));
  XNOR2_X1  g250(.A(new_n352), .B(new_n551), .ZN(new_n552));
  AOI22_X1  g251(.A1(G113), .A2(new_n373), .B1(G5194), .B2(G115), .ZN(new_n553));
  XNOR2_X1  g252(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g253(.A(G130), .B(G132), .ZN(new_n555));
  AOI22_X1  g254(.A1(G117), .A2(new_n388), .B1(new_n393), .B2(G119), .ZN(new_n556));
  XNOR2_X1  g255(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g256(.A(new_n554), .B(new_n557), .Z(new_n558));
  INV_X1    g257(.A(new_n558), .ZN(G5242));
  OAI22_X1  g258(.A1(new_n445), .A2(G90), .B1(G88), .B2(new_n425), .ZN(new_n560));
  XNOR2_X1  g259(.A(G103), .B(new_n560), .ZN(new_n561));
  OAI22_X1  g260(.A1(G92), .A2(G94), .B1(new_n450), .B2(new_n439), .ZN(new_n562));
  XOR2_X1   g261(.A(new_n412), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g262(.A(new_n561), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g263(.A(G109), .B(G111), .ZN(new_n565));
  AOI22_X1  g264(.A1(G105), .A2(new_n431), .B1(new_n399), .B2(G107), .ZN(new_n566));
  XNOR2_X1  g265(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g266(.A(new_n564), .B(new_n567), .Z(G5243));
  OAI22_X1  g267(.A1(G142), .A2(new_n497), .B1(new_n493), .B2(new_n492), .ZN(new_n569));
  NOR2_X1   g268(.A1(new_n411), .A2(new_n470), .ZN(new_n570));
  AOI21_X1  g269(.A(new_n477), .B1(new_n434), .B2(new_n473), .ZN(new_n571));
  NOR2_X1   g270(.A1(new_n466), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g271(.A1(new_n467), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g272(.A1(new_n460), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g273(.A1(new_n462), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g274(.A(new_n471), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  OAI221_X1 g275(.A(new_n569), .B1(new_n444), .B2(new_n496), .C1(new_n508), .C2(new_n576), .ZN(G5244));
  BUF_X1    g276(.A(G5244), .Z(G5246));
  BUF_X1    g277(.A(G5245), .Z(G5247));
  INV_X1    g278(.A(G177), .ZN(new_n580));
  OAI221_X1 g279(.A(G176), .B1(G60), .B2(G177), .C1(new_n580), .C2(new_n369), .ZN(new_n581));
  NOR2_X1   g280(.A1(G176), .A2(new_n580), .ZN(new_n582));
  INV_X1    g281(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g282(.A(G21), .B(new_n534), .ZN(new_n584));
  OAI21_X1  g283(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g284(.A(new_n585), .ZN(G5248));
  OAI221_X1 g285(.A(G176), .B1(G58), .B2(G177), .C1(new_n580), .C2(new_n385), .ZN(new_n587));
  OAI21_X1  g286(.A(new_n533), .B1(G150), .B2(new_n535), .ZN(new_n588));
  XOR2_X1   g287(.A(new_n534), .B(new_n588), .Z(new_n589));
  INV_X1    g288(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g289(.A(new_n587), .B1(new_n583), .B2(new_n590), .ZN(new_n591));
  INV_X1    g290(.A(new_n591), .ZN(G5249));
  OAI221_X1 g291(.A(G176), .B1(G48), .B2(G177), .C1(new_n580), .C2(new_n423), .ZN(new_n593));
  AOI21_X1  g292(.A(new_n476), .B1(new_n421), .B2(new_n475), .ZN(new_n594));
  XNOR2_X1  g293(.A(G2), .B(new_n594), .ZN(new_n595));
  OAI21_X1  g294(.A(new_n593), .B1(new_n583), .B2(new_n595), .ZN(new_n596));
  INV_X1    g295(.A(new_n596), .ZN(G5250));
  INV_X1    g296(.A(G172), .ZN(new_n598));
  INV_X1    g297(.A(G173), .ZN(new_n599));
  OAI221_X1 g298(.A(new_n598), .B1(G22), .B2(G173), .C1(G3), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g299(.A1(G172), .A2(G173), .ZN(new_n601));
  NAND2_X1  g300(.A1(G172), .A2(new_n599), .ZN(new_n602));
  OAI221_X1 g301(.A(new_n600), .B1(G5248), .B2(new_n601), .C1(G5250), .C2(new_n602), .ZN(G5252));
  OAI221_X1 g302(.A(G176), .B1(G19), .B2(G177), .C1(new_n580), .C2(new_n359), .ZN(new_n604));
  INV_X1    g303(.A(new_n604), .ZN(new_n605));
  INV_X1    g304(.A(new_n539), .ZN(new_n606));
  OAI21_X1  g305(.A(new_n538), .B1(G148), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g306(.A(new_n607), .B1(new_n370), .B2(new_n539), .ZN(new_n608));
  NAND2_X1  g307(.A1(new_n544), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g308(.A(new_n609), .B1(new_n544), .B2(new_n608), .ZN(new_n610));
  AOI21_X1  g309(.A(new_n605), .B1(new_n582), .B2(new_n610), .ZN(G5253));
  OAI221_X1 g310(.A(G176), .B1(G59), .B2(G177), .C1(new_n580), .C2(new_n372), .ZN(new_n612));
  INV_X1    g311(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g312(.A(new_n542), .B1(new_n538), .B2(new_n541), .ZN(new_n614));
  AOI21_X1  g313(.A(new_n613), .B1(new_n582), .B2(new_n614), .ZN(G5254));
  OAI221_X1 g314(.A(G176), .B1(G50), .B2(G177), .C1(new_n580), .C2(new_n365), .ZN(new_n616));
  XOR2_X1   g315(.A(new_n530), .B(new_n537), .Z(new_n617));
  OAI21_X1  g316(.A(new_n616), .B1(new_n583), .B2(new_n617), .ZN(new_n618));
  INV_X1    g317(.A(new_n618), .ZN(G5255));
  INV_X1    g318(.A(G175), .ZN(new_n620));
  INV_X1    g319(.A(G174), .ZN(new_n621));
  OAI221_X1 g320(.A(new_n620), .B1(G22), .B2(G174), .C1(G3), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g321(.A1(G174), .A2(G175), .ZN(new_n623));
  NAND2_X1  g322(.A1(new_n621), .A2(G175), .ZN(new_n624));
  OAI221_X1 g323(.A(new_n622), .B1(G5248), .B2(new_n623), .C1(G5250), .C2(new_n624), .ZN(G5256));
  NAND3_X1  g324(.A1(G53), .A2(G176), .A3(new_n580), .ZN(new_n626));
  INV_X1    g325(.A(G176), .ZN(new_n627));
  NOR2_X1   g326(.A1(new_n627), .A2(new_n580), .ZN(new_n628));
  INV_X1    g327(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g328(.A(new_n626), .B1(new_n416), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g329(.A(new_n476), .B1(G2), .B2(new_n594), .ZN(new_n631));
  OAI22_X1  g330(.A1(new_n434), .A2(new_n473), .B1(new_n474), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g331(.A(new_n466), .B1(new_n468), .B2(new_n632), .ZN(new_n633));
  OAI22_X1  g332(.A1(new_n462), .A2(new_n574), .B1(new_n464), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g333(.A1(new_n472), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g334(.A(new_n635), .B1(new_n472), .B2(new_n634), .ZN(new_n636));
  AOI21_X1  g335(.A(new_n630), .B1(new_n582), .B2(new_n636), .ZN(G5257));
  OAI221_X1 g336(.A(G176), .B1(G57), .B2(G177), .C1(new_n580), .C2(new_n410), .ZN(new_n638));
  XOR2_X1   g337(.A(new_n464), .B(new_n633), .Z(new_n639));
  OAI21_X1  g338(.A(new_n638), .B1(new_n583), .B2(new_n639), .ZN(new_n640));
  INV_X1    g339(.A(new_n640), .ZN(G5258));
  OAI221_X1 g340(.A(G176), .B1(G56), .B2(G177), .C1(new_n580), .C2(new_n404), .ZN(new_n642));
  XOR2_X1   g341(.A(new_n468), .B(new_n632), .Z(new_n643));
  OAI21_X1  g342(.A(new_n642), .B1(new_n583), .B2(new_n643), .ZN(new_n644));
  INV_X1    g343(.A(new_n644), .ZN(G5259));
  OAI221_X1 g344(.A(G176), .B1(G55), .B2(G177), .C1(new_n580), .C2(new_n436), .ZN(new_n646));
  XOR2_X1   g345(.A(new_n474), .B(new_n631), .Z(new_n647));
  OAI21_X1  g346(.A(new_n646), .B1(new_n583), .B2(new_n647), .ZN(new_n648));
  INV_X1    g347(.A(new_n648), .ZN(G5260));
  XOR2_X1   g348(.A(G5251), .B(new_n517), .Z(new_n650));
  XNOR2_X1  g349(.A(new_n519), .B(new_n650), .ZN(new_n651));
  OAI22_X1  g350(.A1(new_n510), .A2(G132), .B1(G123), .B2(G133), .ZN(new_n652));
  XNOR2_X1  g351(.A(new_n534), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g352(.A(new_n527), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g353(.A(new_n531), .B(new_n654), .ZN(new_n655));
  OAI22_X1  g354(.A1(new_n539), .A2(new_n543), .B1(G122), .B2(new_n606), .ZN(new_n656));
  XOR2_X1   g355(.A(new_n655), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g356(.A(new_n651), .B(new_n657), .ZN(G5261));
  OAI22_X1  g357(.A1(new_n459), .A2(new_n490), .B1(new_n461), .B2(new_n489), .ZN(new_n659));
  OAI22_X1  g358(.A1(new_n475), .A2(new_n485), .B1(new_n478), .B2(new_n482), .ZN(new_n660));
  XOR2_X1   g359(.A(new_n659), .B(new_n660), .Z(new_n661));
  XNOR2_X1  g360(.A(new_n465), .B(new_n661), .ZN(new_n662));
  AOI22_X1  g361(.A1(G112), .A2(new_n458), .B1(G111), .B2(G124), .ZN(new_n663));
  XNOR2_X1  g362(.A(new_n470), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g363(.A(new_n483), .B(new_n497), .ZN(new_n665));
  XOR2_X1   g364(.A(new_n664), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g365(.A(new_n473), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g366(.A(new_n662), .B(new_n667), .Z(G5262));
  AOI21_X1  g367(.A(new_n635), .B1(new_n411), .B2(new_n470), .ZN(new_n669));
  AOI21_X1  g368(.A(new_n487), .B1(new_n501), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g369(.A1(new_n494), .A2(new_n506), .ZN(new_n671));
  XOR2_X1   g370(.A(new_n670), .B(new_n671), .Z(new_n672));
  NAND4_X1  g371(.A1(new_n595), .A2(new_n647), .A3(new_n643), .A4(new_n639), .ZN(new_n673));
  XNOR2_X1  g372(.A(new_n500), .B(new_n669), .ZN(new_n674));
  NOR3_X1   g373(.A1(new_n636), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g374(.A(new_n669), .ZN(new_n676));
  OAI22_X1  g375(.A1(new_n499), .A2(new_n676), .B1(new_n484), .B2(new_n669), .ZN(new_n677));
  XOR2_X1   g376(.A(new_n486), .B(new_n677), .Z(new_n678));
  AOI21_X1  g377(.A(new_n491), .B1(new_n494), .B2(new_n670), .ZN(new_n679));
  XNOR2_X1  g378(.A(new_n498), .B(new_n679), .ZN(new_n680));
  AND4_X1   g379(.A1(new_n672), .A2(new_n675), .A3(new_n678), .A4(new_n680), .ZN(G5263));
  NOR2_X1   g380(.A1(new_n518), .A2(new_n521), .ZN(new_n682));
  OAI21_X1  g381(.A(new_n609), .B1(new_n356), .B2(new_n543), .ZN(new_n683));
  XNOR2_X1  g382(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND4_X1  g383(.A1(G5251), .A2(new_n584), .A3(new_n590), .A4(new_n617), .ZN(new_n685));
  NOR3_X1   g384(.A1(new_n614), .A2(new_n685), .A3(new_n610), .ZN(new_n686));
  INV_X1    g385(.A(new_n683), .ZN(new_n687));
  NOR2_X1   g386(.A1(new_n518), .A2(new_n687), .ZN(new_n688));
  INV_X1    g387(.A(new_n521), .ZN(new_n689));
  AOI21_X1  g388(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g389(.A(new_n545), .B(new_n690), .ZN(new_n691));
  NOR3_X1   g390(.A1(new_n521), .A2(new_n522), .A3(new_n688), .ZN(new_n692));
  NOR2_X1   g391(.A1(new_n520), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g392(.A(new_n512), .B(new_n693), .Z(new_n694));
  AND4_X1   g393(.A1(new_n684), .A2(new_n686), .A3(new_n691), .A4(new_n694), .ZN(G5264));
  INV_X1    g394(.A(G159), .ZN(new_n696));
  INV_X1    g395(.A(G158), .ZN(new_n697));
  OAI221_X1 g396(.A(new_n696), .B1(G81), .B2(G158), .C1(G80), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g397(.A1(G158), .A2(G159), .ZN(new_n699));
  NAND2_X1  g398(.A1(new_n697), .A2(G159), .ZN(new_n700));
  OAI221_X1 g399(.A(new_n698), .B1(G5248), .B2(new_n699), .C1(G5250), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g400(.A1(G64), .A2(new_n701), .ZN(G5265));
  INV_X1    g401(.A(G161), .ZN(new_n703));
  INV_X1    g402(.A(G160), .ZN(new_n704));
  OAI221_X1 g403(.A(new_n703), .B1(G81), .B2(G160), .C1(G80), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g404(.A1(G160), .A2(G161), .ZN(new_n706));
  NAND2_X1  g405(.A1(new_n704), .A2(G161), .ZN(new_n707));
  OAI221_X1 g406(.A(new_n705), .B1(G5248), .B2(new_n706), .C1(G5250), .C2(new_n707), .ZN(new_n708));
  AND2_X1   g407(.A1(G64), .A2(new_n708), .ZN(G5266));
  OAI221_X1 g408(.A(new_n598), .B1(G14), .B2(G173), .C1(G16), .C2(new_n599), .ZN(new_n710));
  OAI221_X1 g409(.A(new_n710), .B1(new_n601), .B2(G5253), .C1(new_n602), .C2(G5257), .ZN(G5267));
  OAI221_X1 g410(.A(new_n598), .B1(G6), .B2(G173), .C1(G27), .C2(new_n599), .ZN(new_n712));
  OAI221_X1 g411(.A(new_n712), .B1(new_n601), .B2(G5254), .C1(new_n602), .C2(G5258), .ZN(G5268));
  OAI221_X1 g412(.A(new_n598), .B1(G5), .B2(G173), .C1(G26), .C2(new_n599), .ZN(new_n714));
  OAI221_X1 g413(.A(new_n714), .B1(new_n601), .B2(G5255), .C1(new_n602), .C2(G5259), .ZN(G5269));
  OAI221_X1 g414(.A(new_n598), .B1(G25), .B2(G173), .C1(G24), .C2(new_n599), .ZN(new_n716));
  OAI221_X1 g415(.A(new_n716), .B1(G5249), .B2(new_n601), .C1(new_n602), .C2(G5260), .ZN(G5270));
  OAI221_X1 g416(.A(new_n620), .B1(G14), .B2(G174), .C1(G16), .C2(new_n621), .ZN(new_n718));
  OAI221_X1 g417(.A(new_n718), .B1(G5253), .B2(new_n623), .C1(new_n624), .C2(G5257), .ZN(G5271));
  OAI221_X1 g418(.A(new_n620), .B1(G6), .B2(G174), .C1(G27), .C2(new_n621), .ZN(new_n720));
  OAI221_X1 g419(.A(new_n720), .B1(G5254), .B2(new_n623), .C1(new_n624), .C2(G5258), .ZN(G5272));
  OAI221_X1 g420(.A(new_n620), .B1(G5), .B2(G174), .C1(G26), .C2(new_n621), .ZN(new_n722));
  OAI221_X1 g421(.A(new_n722), .B1(G5255), .B2(new_n623), .C1(new_n624), .C2(G5259), .ZN(G5273));
  OAI221_X1 g422(.A(new_n620), .B1(G25), .B2(G174), .C1(G24), .C2(new_n621), .ZN(new_n724));
  OAI221_X1 g423(.A(new_n724), .B1(G5249), .B2(new_n623), .C1(new_n624), .C2(G5260), .ZN(G5274));
  OAI221_X1 g424(.A(new_n696), .B1(G76), .B2(G158), .C1(G86), .C2(new_n697), .ZN(new_n726));
  OAI221_X1 g425(.A(new_n726), .B1(G5253), .B2(new_n699), .C1(G5257), .C2(new_n700), .ZN(new_n727));
  AND2_X1   g426(.A1(G64), .A2(new_n727), .ZN(G5275));
  OAI221_X1 g427(.A(new_n696), .B1(G72), .B2(G158), .C1(G82), .C2(new_n697), .ZN(new_n729));
  OAI221_X1 g428(.A(new_n729), .B1(G5249), .B2(new_n699), .C1(G5260), .C2(new_n700), .ZN(new_n730));
  AND2_X1   g429(.A1(G64), .A2(new_n730), .ZN(G5276));
  OAI221_X1 g430(.A(new_n696), .B1(G70), .B2(G158), .C1(G71), .C2(new_n697), .ZN(new_n732));
  OAI221_X1 g431(.A(new_n732), .B1(G5255), .B2(new_n699), .C1(G5259), .C2(new_n700), .ZN(new_n733));
  AND2_X1   g432(.A1(G64), .A2(new_n733), .ZN(G5277));
  OAI221_X1 g433(.A(new_n696), .B1(G68), .B2(G158), .C1(G69), .C2(new_n697), .ZN(new_n735));
  OAI221_X1 g434(.A(new_n735), .B1(G5254), .B2(new_n699), .C1(G5258), .C2(new_n700), .ZN(new_n736));
  AND2_X1   g435(.A1(G64), .A2(new_n736), .ZN(G5278));
  OAI221_X1 g436(.A(new_n703), .B1(G76), .B2(G160), .C1(G86), .C2(new_n704), .ZN(new_n738));
  OAI221_X1 g437(.A(new_n738), .B1(G5253), .B2(new_n706), .C1(G5257), .C2(new_n707), .ZN(new_n739));
  AND2_X1   g438(.A1(G64), .A2(new_n739), .ZN(G5279));
  OAI221_X1 g439(.A(new_n703), .B1(G72), .B2(G160), .C1(G82), .C2(new_n704), .ZN(new_n741));
  OAI221_X1 g440(.A(new_n741), .B1(G5249), .B2(new_n706), .C1(G5260), .C2(new_n707), .ZN(new_n742));
  AND2_X1   g441(.A1(G64), .A2(new_n742), .ZN(G5280));
  OAI221_X1 g442(.A(new_n703), .B1(G70), .B2(G160), .C1(G71), .C2(new_n704), .ZN(new_n744));
  OAI221_X1 g443(.A(new_n744), .B1(G5255), .B2(new_n706), .C1(G5259), .C2(new_n707), .ZN(new_n745));
  AND2_X1   g444(.A1(G64), .A2(new_n745), .ZN(G5281));
  OAI221_X1 g445(.A(new_n703), .B1(G68), .B2(G160), .C1(G69), .C2(new_n704), .ZN(new_n747));
  OAI221_X1 g446(.A(new_n747), .B1(G5254), .B2(new_n706), .C1(G5258), .C2(new_n707), .ZN(new_n748));
  AND2_X1   g447(.A1(G64), .A2(new_n748), .ZN(G5282));
  INV_X1    g448(.A(G170), .ZN(new_n750));
  AOI221_X1 g449(.A(G171), .B1(G54), .B2(G170), .C1(new_n750), .C2(new_n378), .ZN(new_n751));
  XOR2_X1   g450(.A(G61), .B(new_n511), .Z(new_n752));
  OAI221_X1 g451(.A(G171), .B1(new_n750), .B2(G5251), .C1(G170), .C2(new_n752), .ZN(new_n753));
  INV_X1    g452(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g453(.A(new_n751), .B(new_n754), .C1(G62), .C2(G178), .ZN(G5283));
  XOR2_X1   g454(.A(G61), .B(new_n512), .Z(G5284));
  OAI221_X1 g455(.A(G176), .B1(G54), .B2(G177), .C1(new_n580), .C2(new_n378), .ZN(new_n757));
  OAI21_X1  g456(.A(new_n757), .B1(G5251), .B2(new_n583), .ZN(new_n758));
  INV_X1    g457(.A(new_n758), .ZN(G5285));
  OAI221_X1 g458(.A(G176), .B1(G52), .B2(G177), .C1(new_n580), .C2(new_n374), .ZN(new_n760));
  OAI21_X1  g459(.A(new_n760), .B1(new_n583), .B2(new_n694), .ZN(new_n761));
  INV_X1    g460(.A(new_n761), .ZN(G5286));
  OAI221_X1 g461(.A(G176), .B1(G47), .B2(G177), .C1(new_n580), .C2(new_n396), .ZN(new_n763));
  OAI21_X1  g462(.A(new_n763), .B1(new_n583), .B2(new_n691), .ZN(new_n764));
  INV_X1    g463(.A(new_n764), .ZN(G5287));
  OAI221_X1 g464(.A(G176), .B1(G43), .B2(G177), .C1(new_n580), .C2(new_n391), .ZN(new_n766));
  OAI21_X1  g465(.A(new_n766), .B1(new_n583), .B2(new_n684), .ZN(new_n767));
  INV_X1    g466(.A(new_n767), .ZN(G5288));
  NAND3_X1  g467(.A1(G99), .A2(G155), .A3(G5199), .ZN(new_n769));
  NOR3_X1   g468(.A1(G5213), .A2(new_n769), .A3(new_n558), .ZN(new_n770));
  AND4_X1   g469(.A1(G5243), .A2(new_n770), .A3(G5262), .A4(G5261), .ZN(G5289));
  INV_X1    g470(.A(new_n448), .ZN(new_n772));
  OAI221_X1 g471(.A(G176), .B1(G46), .B2(G177), .C1(new_n580), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g472(.A(new_n773), .B1(new_n583), .B2(new_n680), .ZN(new_n774));
  INV_X1    g473(.A(new_n774), .ZN(G5290));
  NAND3_X1  g474(.A1(G45), .A2(G176), .A3(new_n580), .ZN(new_n776));
  OAI221_X1 g475(.A(new_n776), .B1(new_n429), .B2(new_n629), .C1(new_n583), .C2(new_n672), .ZN(new_n777));
  INV_X1    g476(.A(new_n777), .ZN(G5291));
  NAND3_X1  g477(.A1(G20), .A2(G176), .A3(new_n580), .ZN(new_n779));
  OAI221_X1 g478(.A(new_n779), .B1(new_n454), .B2(new_n629), .C1(new_n583), .C2(new_n678), .ZN(new_n780));
  INV_X1    g479(.A(new_n780), .ZN(G5292));
  NAND3_X1  g480(.A1(G44), .A2(G176), .A3(new_n580), .ZN(new_n782));
  OAI21_X1  g481(.A(new_n782), .B1(new_n443), .B2(new_n629), .ZN(new_n783));
  AOI21_X1  g482(.A(new_n783), .B1(new_n582), .B2(new_n674), .ZN(G5293));
  OAI221_X1 g483(.A(new_n620), .B1(G41), .B2(G174), .C1(G42), .C2(new_n621), .ZN(new_n785));
  OAI221_X1 g484(.A(new_n785), .B1(new_n623), .B2(G5285), .C1(new_n624), .C2(G5290), .ZN(G5294));
  OAI221_X1 g485(.A(new_n598), .B1(G41), .B2(G173), .C1(G42), .C2(new_n599), .ZN(new_n787));
  OAI221_X1 g486(.A(new_n787), .B1(new_n601), .B2(G5285), .C1(new_n602), .C2(G5290), .ZN(G5295));
  OAI221_X1 g487(.A(new_n598), .B1(G18), .B2(G173), .C1(G17), .C2(new_n599), .ZN(new_n789));
  OAI221_X1 g488(.A(new_n789), .B1(new_n601), .B2(G5286), .C1(new_n602), .C2(G5291), .ZN(G5296));
  OAI221_X1 g489(.A(new_n598), .B1(G40), .B2(G173), .C1(G39), .C2(new_n599), .ZN(new_n791));
  OAI221_X1 g490(.A(new_n791), .B1(new_n601), .B2(G5287), .C1(new_n602), .C2(G5292), .ZN(G5297));
  OAI221_X1 g491(.A(new_n598), .B1(G15), .B2(G173), .C1(G36), .C2(new_n599), .ZN(new_n793));
  OAI221_X1 g492(.A(new_n793), .B1(new_n601), .B2(G5288), .C1(new_n602), .C2(G5293), .ZN(G5298));
  OAI221_X1 g493(.A(new_n620), .B1(G18), .B2(G174), .C1(G17), .C2(new_n621), .ZN(new_n795));
  OAI221_X1 g494(.A(new_n795), .B1(new_n623), .B2(G5286), .C1(new_n624), .C2(G5291), .ZN(G5299));
  OAI221_X1 g495(.A(new_n620), .B1(G40), .B2(G174), .C1(G39), .C2(new_n621), .ZN(new_n797));
  OAI221_X1 g496(.A(new_n797), .B1(new_n623), .B2(G5287), .C1(new_n624), .C2(G5292), .ZN(G5300));
  OAI221_X1 g497(.A(new_n620), .B1(G15), .B2(G174), .C1(G36), .C2(new_n621), .ZN(new_n799));
  OAI221_X1 g498(.A(new_n799), .B1(new_n623), .B2(G5288), .C1(new_n624), .C2(G5293), .ZN(G5301));
  OAI221_X1 g499(.A(new_n696), .B1(G77), .B2(G158), .C1(G87), .C2(new_n697), .ZN(new_n801));
  OAI221_X1 g500(.A(new_n801), .B1(new_n699), .B2(G5288), .C1(new_n700), .C2(G5293), .ZN(new_n802));
  AND2_X1   g501(.A1(G64), .A2(new_n802), .ZN(G5302));
  OAI221_X1 g502(.A(new_n696), .B1(G75), .B2(G158), .C1(G85), .C2(new_n697), .ZN(new_n804));
  OAI221_X1 g503(.A(new_n804), .B1(new_n699), .B2(G5287), .C1(new_n700), .C2(G5292), .ZN(new_n805));
  AND2_X1   g504(.A1(G64), .A2(new_n805), .ZN(G5303));
  OAI221_X1 g505(.A(new_n696), .B1(G74), .B2(G158), .C1(G84), .C2(new_n697), .ZN(new_n807));
  OAI221_X1 g506(.A(new_n807), .B1(new_n699), .B2(G5286), .C1(new_n700), .C2(G5291), .ZN(new_n808));
  AND2_X1   g507(.A1(G64), .A2(new_n808), .ZN(G5304));
  OAI221_X1 g508(.A(new_n696), .B1(G73), .B2(G158), .C1(G83), .C2(new_n697), .ZN(new_n810));
  OAI221_X1 g509(.A(new_n810), .B1(new_n699), .B2(G5285), .C1(new_n700), .C2(G5290), .ZN(new_n811));
  AND2_X1   g510(.A1(G64), .A2(new_n811), .ZN(G5305));
  OAI221_X1 g511(.A(new_n703), .B1(G77), .B2(G160), .C1(G87), .C2(new_n704), .ZN(new_n813));
  OAI221_X1 g512(.A(new_n813), .B1(new_n706), .B2(G5288), .C1(new_n707), .C2(G5293), .ZN(new_n814));
  AND2_X1   g513(.A1(G64), .A2(new_n814), .ZN(G5306));
  OAI221_X1 g514(.A(new_n703), .B1(G75), .B2(G160), .C1(G85), .C2(new_n704), .ZN(new_n816));
  OAI221_X1 g515(.A(new_n816), .B1(new_n706), .B2(G5287), .C1(new_n707), .C2(G5292), .ZN(new_n817));
  AND2_X1   g516(.A1(G64), .A2(new_n817), .ZN(G5307));
  OAI221_X1 g517(.A(new_n703), .B1(G74), .B2(G160), .C1(G84), .C2(new_n704), .ZN(new_n819));
  OAI221_X1 g518(.A(new_n819), .B1(new_n706), .B2(G5286), .C1(new_n707), .C2(G5291), .ZN(new_n820));
  AND2_X1   g519(.A1(G64), .A2(new_n820), .ZN(G5308));
  OAI221_X1 g520(.A(new_n703), .B1(G73), .B2(G160), .C1(G83), .C2(new_n704), .ZN(new_n822));
  OAI221_X1 g521(.A(new_n822), .B1(new_n706), .B2(G5285), .C1(new_n707), .C2(G5290), .ZN(new_n823));
  AND2_X1   g522(.A1(G64), .A2(new_n823), .ZN(G5309));
  AOI222_X1 g523(.A1(new_n521), .A2(new_n523), .B1(new_n689), .B2(new_n522), .C1(new_n518), .C2(new_n545), .ZN(new_n825));
  XNOR2_X1  g524(.A(new_n511), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g525(.A(G5251), .B(new_n526), .ZN(new_n827));
  OAI22_X1  g526(.A1(new_n687), .A2(new_n826), .B1(new_n683), .B2(new_n827), .ZN(new_n828));
  INV_X1    g527(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g528(.A(new_n607), .B1(new_n538), .B2(new_n540), .ZN(new_n830));
  INV_X1    g529(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g530(.A(new_n536), .B1(new_n532), .B2(new_n534), .ZN(new_n832));
  XOR2_X1   g531(.A(new_n831), .B(new_n832), .Z(new_n833));
  INV_X1    g532(.A(new_n833), .ZN(new_n834));
  AOI221_X1 g533(.A(G162), .B1(new_n589), .B2(new_n833), .C1(new_n590), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g534(.A(G162), .B1(new_n588), .B2(new_n831), .ZN(new_n836));
  AOI21_X1  g535(.A(new_n836), .B1(new_n588), .B2(new_n834), .ZN(new_n837));
  NOR2_X1   g536(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g537(.A(new_n530), .B(new_n838), .Z(new_n839));
  XOR2_X1   g538(.A(new_n544), .B(new_n839), .Z(new_n840));
  XNOR2_X1  g539(.A(new_n541), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g540(.A(new_n582), .B1(new_n829), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g541(.A(new_n842), .B1(new_n829), .B2(new_n841), .ZN(new_n843));
  XNOR2_X1  g542(.A(new_n391), .B(new_n396), .ZN(new_n844));
  OAI21_X1  g543(.A(new_n379), .B1(new_n375), .B2(new_n378), .ZN(new_n845));
  XNOR2_X1  g544(.A(new_n844), .B(new_n845), .ZN(new_n846));
  OAI22_X1  g545(.A1(G100), .A2(new_n370), .B1(new_n377), .B2(G148), .ZN(new_n847));
  AOI221_X1 g546(.A(new_n356), .B1(new_n368), .B2(new_n352), .C1(new_n366), .C2(G121), .ZN(new_n848));
  AOI221_X1 g547(.A(G147), .B1(G98), .B2(new_n352), .C1(G102), .C2(G121), .ZN(new_n849));
  OR2_X1    g548(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI221_X1 g549(.A(new_n363), .B1(new_n368), .B2(new_n360), .C1(new_n366), .C2(G126), .ZN(new_n851));
  AOI221_X1 g550(.A(G149), .B1(G98), .B2(new_n360), .C1(G102), .C2(G126), .ZN(new_n852));
  OR2_X1    g551(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI221_X1 g552(.A(new_n383), .B1(new_n368), .B2(new_n380), .C1(new_n366), .C2(G128), .ZN(new_n854));
  AOI221_X1 g553(.A(G150), .B1(G98), .B2(new_n380), .C1(G102), .C2(G128), .ZN(new_n855));
  NOR2_X1   g554(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g555(.A(new_n369), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g556(.A(new_n853), .B(new_n857), .Z(new_n858));
  XNOR2_X1  g557(.A(new_n850), .B(new_n858), .ZN(new_n859));
  XOR2_X1   g558(.A(new_n847), .B(new_n859), .Z(new_n860));
  OAI21_X1  g559(.A(new_n628), .B1(new_n846), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g560(.A(new_n861), .B1(new_n846), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g561(.A1(new_n843), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g562(.A1(G51), .A2(new_n627), .ZN(new_n864));
  OAI21_X1  g563(.A(new_n863), .B1(G177), .B2(new_n864), .ZN(G5310));
  INV_X1    g564(.A(G157), .ZN(new_n866));
  OAI21_X1  g565(.A(new_n576), .B1(new_n866), .B2(new_n481), .ZN(new_n867));
  INV_X1    g566(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g567(.A(new_n507), .B1(new_n495), .B2(new_n501), .ZN(new_n869));
  XNOR2_X1  g568(.A(new_n498), .B(new_n502), .ZN(new_n870));
  XNOR2_X1  g569(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g570(.A(new_n495), .B(new_n505), .ZN(new_n872));
  OAI22_X1  g571(.A1(new_n868), .A2(new_n871), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g572(.A(new_n467), .B1(new_n479), .B2(new_n572), .ZN(new_n874));
  INV_X1    g573(.A(new_n874), .ZN(new_n875));
  OAI33_X1  g574(.A1(new_n408), .A2(new_n459), .A3(new_n874), .B1(G137), .B2(new_n461), .B3(new_n875), .ZN(new_n876));
  AOI21_X1  g575(.A(new_n477), .B1(new_n474), .B2(new_n476), .ZN(new_n877));
  INV_X1    g576(.A(new_n479), .ZN(new_n878));
  XNOR2_X1  g577(.A(new_n472), .B(new_n571), .ZN(new_n879));
  OAI21_X1  g578(.A(new_n480), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g579(.A(new_n877), .B(new_n880), .ZN(new_n881));
  XOR2_X1   g580(.A(new_n876), .B(new_n881), .Z(new_n882));
  INV_X1    g581(.A(new_n594), .ZN(new_n883));
  AOI21_X1  g582(.A(new_n878), .B1(new_n883), .B2(new_n877), .ZN(new_n884));
  INV_X1    g583(.A(new_n462), .ZN(new_n885));
  AOI21_X1  g584(.A(new_n574), .B1(new_n885), .B2(new_n573), .ZN(new_n886));
  XNOR2_X1  g585(.A(new_n879), .B(new_n886), .ZN(new_n887));
  XOR2_X1   g586(.A(new_n884), .B(new_n887), .Z(new_n888));
  OAI22_X1  g587(.A1(new_n866), .A2(new_n882), .B1(G157), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g588(.A1(new_n463), .A2(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n890));
  XNOR2_X1  g589(.A(new_n671), .B(new_n890), .ZN(new_n891));
  XOR2_X1   g590(.A(new_n889), .B(new_n891), .Z(new_n892));
  NOR2_X1   g591(.A1(new_n873), .A2(new_n892), .ZN(new_n893));
  AOI211_X1 g592(.A(new_n583), .B(new_n893), .C1(new_n873), .C2(new_n892), .ZN(new_n894));
  OAI221_X1 g593(.A(new_n438), .B1(G94), .B2(G98), .C1(new_n439), .C2(G102), .ZN(new_n895));
  OAI221_X1 g594(.A(new_n895), .B1(G100), .B2(new_n441), .C1(G101), .C2(new_n442), .ZN(new_n896));
  XNOR2_X1  g595(.A(new_n448), .B(new_n896), .ZN(new_n897));
  OAI221_X1 g596(.A(new_n424), .B1(G90), .B2(G98), .C1(new_n425), .C2(G102), .ZN(new_n898));
  OAI221_X1 g597(.A(new_n898), .B1(G100), .B2(new_n427), .C1(G101), .C2(new_n428), .ZN(new_n899));
  OAI221_X1 g598(.A(new_n449), .B1(G92), .B2(G98), .C1(new_n450), .C2(G102), .ZN(new_n900));
  OAI221_X1 g599(.A(new_n900), .B1(G100), .B2(new_n452), .C1(G101), .C2(new_n453), .ZN(new_n901));
  XOR2_X1   g600(.A(new_n899), .B(new_n901), .Z(new_n902));
  XOR2_X1   g601(.A(new_n897), .B(new_n902), .Z(new_n903));
  AOI221_X1 g602(.A(new_n434), .B1(new_n368), .B2(new_n431), .C1(new_n366), .C2(G107), .ZN(new_n904));
  AOI221_X1 g603(.A(G139), .B1(G98), .B2(new_n431), .C1(G102), .C2(G107), .ZN(new_n905));
  NOR2_X1   g604(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI221_X1 g605(.A(new_n402), .B1(new_n368), .B2(new_n399), .C1(new_n366), .C2(G105), .ZN(new_n907));
  AOI221_X1 g606(.A(G138), .B1(G98), .B2(new_n399), .C1(G102), .C2(G105), .ZN(new_n908));
  OR2_X1    g607(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g608(.A(new_n906), .B(new_n909), .ZN(new_n910));
  AOI221_X1 g609(.A(new_n408), .B1(new_n368), .B2(new_n405), .C1(new_n366), .C2(G103), .ZN(new_n911));
  AOI221_X1 g610(.A(G137), .B1(G98), .B2(new_n405), .C1(G102), .C2(G103), .ZN(new_n912));
  NOR2_X1   g611(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g612(.A(new_n910), .B(new_n913), .ZN(new_n914));
  AOI221_X1 g613(.A(new_n421), .B1(new_n368), .B2(new_n418), .C1(new_n366), .C2(G109), .ZN(new_n915));
  AOI221_X1 g614(.A(G135), .B1(G98), .B2(new_n418), .C1(G102), .C2(G109), .ZN(new_n916));
  OR2_X1    g615(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI221_X1 g616(.A(new_n411), .B1(G96), .B2(G98), .C1(new_n412), .C2(G102), .ZN(new_n918));
  OAI221_X1 g617(.A(new_n918), .B1(G100), .B2(new_n414), .C1(G101), .C2(new_n415), .ZN(new_n919));
  XOR2_X1   g618(.A(new_n917), .B(new_n919), .Z(new_n920));
  XOR2_X1   g619(.A(new_n914), .B(new_n920), .Z(new_n921));
  NOR2_X1   g620(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  AOI211_X1 g621(.A(new_n629), .B(new_n922), .C1(new_n903), .C2(new_n921), .ZN(new_n923));
  NOR2_X1   g622(.A1(new_n894), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g623(.A1(G49), .A2(new_n627), .ZN(new_n925));
  OAI21_X1  g624(.A(new_n924), .B1(G177), .B2(new_n925), .ZN(G5311));
  OAI221_X1 g625(.A(new_n598), .B1(G23), .B2(G173), .C1(G4), .C2(new_n599), .ZN(new_n927));
  AOI22_X1  g626(.A1(G38), .A2(new_n580), .B1(G177), .B2(new_n924), .ZN(new_n928));
  AOI22_X1  g627(.A1(G37), .A2(new_n580), .B1(G177), .B2(new_n863), .ZN(new_n929));
  OAI221_X1 g628(.A(new_n927), .B1(new_n602), .B2(new_n928), .C1(new_n601), .C2(new_n929), .ZN(G5312));
  OAI221_X1 g629(.A(new_n620), .B1(G23), .B2(G174), .C1(G4), .C2(new_n621), .ZN(new_n931));
  OAI221_X1 g630(.A(new_n931), .B1(new_n624), .B2(new_n928), .C1(new_n623), .C2(new_n929), .ZN(G5313));
  OAI221_X1 g631(.A(new_n696), .B1(G79), .B2(G158), .C1(G78), .C2(new_n697), .ZN(new_n933));
  OAI221_X1 g632(.A(new_n933), .B1(new_n700), .B2(new_n928), .C1(new_n699), .C2(new_n929), .ZN(new_n934));
  NAND2_X1  g633(.A1(G64), .A2(new_n934), .ZN(G5314));
  OAI221_X1 g634(.A(new_n703), .B1(G79), .B2(G160), .C1(G78), .C2(new_n704), .ZN(new_n936));
  OAI221_X1 g635(.A(new_n936), .B1(new_n707), .B2(new_n928), .C1(new_n706), .C2(new_n929), .ZN(new_n937));
  NAND2_X1  g636(.A1(G64), .A2(new_n937), .ZN(G5315));
endmodule


